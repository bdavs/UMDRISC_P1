XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2���)>�ѱ-�kBd�����D>�T@�<�����Ce$�^i戝��<;YJ6�]5�ﰻ�L��ʦĔ6;��U�eB-h�Rd�/5�*S������(�� ����jF5ɏӺ,�n�,`zM����7����J�9���y�Q���������c]}�o��r��<�Gu����@+@�����8o;�s���LI�I�U�T����L��E%��f�3�:ԋ�Ve�kZd[�Ū9�=Z���ԃ�*-r���'5����t��(pd�%s7Ol����n��O8�Q�2pd��V֯i��3��X%�q�cn�
�,����q;�N�56��Ъ����DB{���� b��1��ė0$�&0H�U�u�i_y������fmFI����e�ò]�5G�LR�0�<�8��QCOZ2�/�ef�éƲ���� �+|��R2�P���T@
�сƝbD(y��k�@��SM�� C_{�#γZQ[�Bk��'oٱ-���!��~ �q�A���ӥf�p�˕"L����9���Iu�1��ު������ծǿ���`�/�$�z�MXH����K�1Z�oub<���J� @ �*�QXT{�KRr&��|h�n$:���\�w��v6��+$�V9H^�̭�ŕB���T�C��[���M,ܟ�P2�t뻺E,��e�R����_ѷ؂��2�}i��	e􅄮 �S�j�C+��X6n���Y�}�E�� �c�B�~R�l)J�G�XlxVHYEB    4089     e40������58���c��/^@U��>ǂ~�9��	���rLxЛ%���B�l�I���~��0�F�/��:�>~�mRO|jS?�x1���2���b����_ 00g�ۢO�g�
�1�"Ǫ#Mۛ�\�Z���n��w=4M9����w/쉎U�6lb����-�O�x�����*e��g}f�>����#����N�IZT�C�$��O��\.�U��Y	07 v��"�Sp�;e����*�Ƥ�z�K��D�� ?u�Po�f��u�V}�?�8���_;!��.�`'GT���ʐ�Hϑ��T�͋|Qq�W��X�����R\J�=[��ϡ��q�p�x�,M_��^�F�R#mQ���Y�rW"+��h�U�x�rv���U�@���U0c�	aE�b(�Ҵ�~�5�{ k�)���O�����*"�����gY��O\zj�0v�T���R�H������C!05������ra�[q/څ�_^���2���iF�q�x��&�(�W���O����!������2>���6 PX�&1a��2`u�~��$�����.�l�A�.�^�H���d����_�>+�7��.v%�&�_�v�%��f�����	�XV���~(z��1Q���u��d�����⚜�>-����q�JZ���v�Ÿ�g�w��
�Z��j^o/�w����e�����Qs�d�ͻ���LK�_�CӔ
Ƣ���{�B֍�!b
^E��5DCI�~�y���I���oCKC�v�}�eBO��I�㇀k��S�rfcGG�yI�Ԝ�T�<V�B]1?q7m0��Wog8k*�+m��=����Y[t�BT�p�q�v���]K̪�#H�oP��Wp"�Ft,k�1����?�װ^�X�ٯX �pX��@���}R���U'k�a�P�r����˲�����¬�eXӣ�A�U,�W0(��ǉ5Oɲ:�͠ ����Q�[�`�
J,����"v���ŕ��ʣ��Ӳ�*Y�-���Ra�2�uy�O���nG���sa���9�G���I��u��Y � �u���T��'S6�2��߲�����7� �+�<6u?������6�2<�y� ��1W�dF�L<���桦�N�ϯ�'��_�n�\���9����̐v1��nJ���RT�w�ܸ�{�I��Q9��ln�HUo�ֈ-:�I�́z�`�Ft�JH�Xi��[>���T���vͱw�7��ȍ�x�����]/qQ���n�?L�0��s���Қ���%=4�{$vBXZ�#���~|b�q�i�GiV.�I-	j���I����*˰ԥ5�U&V8�@/�p��^#Z��+�-W���c��rC��h���o����#'�1���?��yM��$L�������sq�3Q��~.��*�?Pn�%�vC�W�����Y}�xV��ᜢ�î�H�o��lh.
�P�ID_!|}UV+�t �W���i{"�i煢S��w����tΧp�Yr-X����_x5��(jgz����zP�L���Zn뉲?�]n�K�0\hCD�{�L����8��U�s����V��V�c�`��.g�7��k0�����������x�����3Q~qO���=U��r8�L:bTn<�;/�_۪}�\Xت��#�.��K=�8�@L�q�s��P��ޑ�\6�ĲX�3�5w]�Z�P;+$� �����b��l�D u�t$h^Է *���"�{1�T���_j�M�Z�Z�����Rb�-��\]���+�Yn�/�:������-��!C�Q"Y'쵾�ѻйp'�E�4l8'���-�{L��Α�����u"8�s����K������V��g����J/T��� h�:�8	c���D���J�Wm�t�5��g���.H��t?��P�=1�j�0��5�h/���H
��.��xr��:t�ڷM4yr�l���-y��{Z-�q*�+(�+	���K*���W涌c�=���Zl��^jNg$D.2ս9�@�܉�DP�4���/i��[��;�`<��q�9+ �<�#��p���I������7��Ӷ��T]MW<�
�G�\�F�f�T��(Q���|Sh�N��e���4m6mn�x��:��N�k���1����y���^35�ج<���
�-|� ? �~\b0Sv{��MwׁU�n��oJI؝��ڨ�D O�!�<)�!y�؂Q�],��XNß��Gֵ�Pk��lZD]OV��'D���o�����>JL1[|7�e�sj��H��s�6�pk寍*�/��*���0@���}p5��g]q%���'̻��~��a�G^)������t2���a11^��yY�REÌ���ߎU�����2�v %(�$��1������Aq��2�k�~VZ'J�r���Z�,��$Cp"��U�G�jt��%�+��ȳ"G��w�)i�gv��v#�7�A[�R�%8�q�t"�u�1�3�҄*l�1�{A!AG�$�z��?�v��3�]20���8`�h.
#Hߍ�,~Ź�B�0��^�Z��Od�2`s�I�i��'J�8SD"[�.�:��uVP�ՙ� 8�!��m��Z��t��Sy 2������N].E��X������g�_x r���Q�Bu4E�����|��y,���F-xQ�+�;��-��c��G2_yF/���Z9@��G3���{Ұ�w�nM�۬�ٰ���ݎ�T
���9�Ҩ��,!ﱒf�����I����&�u�=����G�t4e�mQ�C'���x:��7��B����Z~f*u/=$*rФG
��(�w��"mQC�;8�N՘�F~q��ײ��g����Y��h{|*-��V��@T��Z�\j�ߕ9<� /�`� ��*��}*G�Y�$n�z�=Jf�V�4᷾12�)���A{2�D3�!�y>��I�L`qN�� �����zz��㳙Q�r���{9V�����tu8��߄��}ݨ��My�"]�T5��G'6P� �s��?A)�B���+	�h5c����gZ{��Ef*������b.Z�P�h�|)��
6��1R�i��yǳv�X��I����A&�����Q�*.a��C�@�qu�;��A|L?uaO�ѡ�SY���
/�����b�3�������x.�_���	i��D�9����E2_��Л�et!�X���!��޷
�a�
d��!��' `��AdI���dU�֙��W�_�D�Jސɍ�1<W�U��f6�.6�����!~�,�T�>nѤ$��n�}�i����єgwe���d��ߨo���Mΐ���t�B�^ �����w�ߦ�ƺ��*T(����c�
�KXem+�p;[Me�D#��|Ӕ�'e��aՔ4���d�gKi��0��2<�.���uQ�(Tۭ��ӄ3�}B�/�"fR~� ���݀�f�BE������H�8��bl��Xxl|Њ
�_��� ���S��-c�s�����=�h��Y}:�<�޾�@~�g�Ѹ4�4�~TZ��8��$�iį�[��[<Ą��@�cL3���#m��+�&�;�t�O�1�Su.k