XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z��sdJ�t���q�2�8c"�{������w���۔�чV07��}���8�B�t����|�R�:'���t���G�:����Q�d<��>-'^4uȡi�o�qc~8vs��[��8��S-�����$�:/4]�wҦ�ׂR�����O���3>�
|�00��G��b��������{)�H�dd����Yg^c�u>��Q��D�*
��x�ڒ����P��e|S@��%݇a��e8;��5 �]Ue0	UR��K�.=D�GW�߬��p�w�R���J�D�����<�W�5`��)C�~�<�?�o��f��.�Dnӻ�ͪ  q�w��%%�]�.�,�ɿ�8�P(�p�n������ ��Dib��V�h�RjVt�+]�?ͣ�ܭe��0Sp,I�Z.��i�CPv��9Ǘ�H}��O�C�<�AR�羇5E��|FeѵH5���3ç��C0�F�b����\��v�.��+s�D�����r���J���jk'1U���5KVs��#���L:q���|.t��6A��+?39j�N��e�
��G��'|���s�>ԁ'�dp+�W�i>�f�4%�7G
k��a���xv�Q��`M� ��<X�o���+P��FT��=�KfB�x� U���[�AP1׈��x4Pi5��j�d�ymm�	�`�Q@>�Q��$=_*��l��xa�%����Fɵ=N�H����s�V�l�,����	:��Ge�v�o�닸�_2
Bj��l�5[�eXlxVHYEB    fa00    1790�f����).m����rʢ���@߸��W�*�S��cuX����PŲ
����[�
]3��?������~�ǁ.zm�����RK;��e�cL���ꂰ�a���U½�yݘu�V{%�Ӿ����X-h)4�@хd���B@%�R�/{`"������?F��&�:ӧ���%�2:��_��ZXP����-v"�&8�u�Q�f��k�l�2���I?���J�~���_[��>Rl�c�VM�G�9�O��ŕ{�sm����������L�M���0 zi%{$T�W�w���?dM/��}ΒP�����>�sma�/sb3�&�?�0Yœ�z�"�hK"Ӑz筱 �Q�7g�s�Kȧ�+SU9.���j��+���EN?�%3y��8�p%�gPO����`�ք�{�z�#�FM��_��_tU�N��Zj�� b4\F
�A��!�i V��h�a!��V�� �W�!8�9�T#"q��ce�z�[��}/�G��)�?t�~�dl2XG*���}Աƌ0�vEO��c/�?F?���4p�|~�ٽD����3?f%��7�jW��,�/!D�iq!�'���G<:-��ژ���^�ձ���ᡜ)+Fqf�R*���Ƒ��ʖå�s�߂�Y��sMwZf뿍���Uu"��[���y�D�<k��ٵ|$ƛ��tL����s�Z}���"[U�d���x3�r
y�:�p�"�]�y@vX�ga�3���W��������y�̻�� �`��e��dW,�Wz�I�Z6:g	��(�~z��B����e\:�/��?�{����̙�͉�"�a��Ke��^�N\��k�VS���A'5� ]Hq�
t�����L�?�I�S���>/�&��l�f>���f� �����R�/�)>���Rs*����^?]�V�k�Eȋ����pu�8��h�.�W���n<�z��M3���q�׋�Πc~�4��#c�%,��$��cb�?�����Xޖ�FӀ�ϝ	��N;�����_�d�~s�<06V֌�EXҡ8������Ќf�<h�?7[�@���n�)���C��^h 4m>o�W체�y?S��s��!>X�=�N�No����@��ȁ��
�OL��jB�c�cA�FmQ�ir�n�Đ�1�	����;�Ѫ�?�[Aɧ7QR���}�4�C���$�.%p~Z*��9Y�0��P�Z�7��iۄX��Mq���Ѿ8��t7m��
���O�+����T���~�L���dD(H�cDg��*d�l]��wsA��.x!	^�����^HH�:�r p)�!�L��t��8���:��� !���5�(S�h	����CN ��k���?\����pkM��k�na��^K[;���A��de�C�7K�
8\I\Yz= ���ު��B�����M���'R:'~.�簃�H�'�)��[Y	�8I����U���B���N1ѳ�q"g{*4�"tU,P��{��?������?��z&�0?�P(������7��h%�W� (�!�A�*M��5|�R���J)~m�a��"� �5w'�~b��&�$�QI�ħ��o�PTegR"���]�SR�k����#h+�DL$ޜ���F�@�L���vm�I�[�������g�:#��n�^�$��_��Яr@@�4��.���Ȥk��������D�_��9�p�vn(9��j�����o3��3���fC�7�I|+��p�o9=f��Geʐ���D���p�E��\��*�G�nin��^$�E��{v=i�6�S&z��������Se�����j;:_p��y�ө���_�%��G��ZWi���:S�&�T({ c.�D��t�*���~)�� r�ʵ�h8m�J�+��2[x�{,S�����!^
	�"���M�L��#v�LƯ��$���rx�1v��/�k#}�A���ٔ���a,������3�jQ�@��nf�쒢@z�2Uy@R�uw���Vy�תt�1����Ҝ+��g�@��j]:(��h���:�^~�Jfǉ�}Y��.U��3A�e"x آx(���Tӕ��B �
W5?H��4�������}��ͨz#PdC��1�R��rl5���X�O�|K5;�9�݊��-t�����f����&��H>$�Bw	� >�p@�US��� �Ă��M�V$15h���ԕM�R��[���#'9�/�-�AsfZ(M輄��s2��܌#e2���.Uڜ��Y��v4K���8o�P��k�D��h����E�r�ÔA��P�o�&`��f���=�rp�F�|n3��t�x8��k�/@;�i�SD;i@�}*���֒#<�?=*+��}�H���RF�t����1)8�>�NL��P�U{K%�0�ȋ^���4�xj
jO�P%��(p��4�M�����
y���f��G�J��ieg�3y��f�޻V�������Ct������dO��[�v%��yc*��xRˉ��J�>�KI�C�Si L��α���Գ:3ƒ�V=���l�TyiMQ/�TJ�>��!ҞH���lV�`W�����j�ث��U�U��^�"S^��Q��6�����}�T0�\B��$�s\������1>���Ƥzᕪ�Q�D���y=-�ӵ!�΂`�U�e�q��ve�$���U6s�h�v �*���a�H��P6���3�_��p1���=�yZ_�U�VR<I�dJ��h�/��E�8�.�W���?�suJit[կP`�T�i�;/�$q�n��4}����>;���T�nZ�0�2X�)�mů��K{g��O��7�B"��_Ls����}���Q�����*��yS�Y���m+!Ǖkޑ��Kc���.'|�l���ɀ:��.2}cO�;K�f �f��ش7s��W��d1�I[��������G��F���ӻ▜@���V�
��а�)#&`q��B��u}~��aG���nQ�ݺh���,�a;�'x��h�~���2�j[MTr�S�Ke8ܸ��A�^ׅ}:���w��ӈ����������R�p&�@�Ys&z"kW* [�4�A�<�����gW�!�_�qM4#7�ӌ[)v5l{O�����)�f[�5qj� V5�(M��EtZ'���9qL��áϘ;��Z&*��r{���_(�UN��*������4o��־x��I�1
˄k�{~�wa���!�T�<�� i�M-��'���;n��TR����^�����R#���oK��be���އF���Xk^n�_ �	�ڦ=J}!���_�gD��s�.�i�'V�䃎����1	0�h�fPJ���}�~d��;�Էޯi�r�A�V-�62݂����$!w*Uf�������p-
�W��$ؚ���N��a�V$"l<U]f܁��~�'�M�\_�_r�'|��G���"+��m��Ǽl�i1&_S����^��pQ���h>�&A>�>�%��t�o�57�n��)�H�ʓ�G$�� R����a}��+��H[w�I�*�&�2��ʗ�����=D�Ї#��	=A����Sm��g׿e�/~,g6��Y!���c�5W����c5]{�e��睩�p����h��(��ppu�Vӹ6�g`� �P,���(�颖?w�`�I�Ζ�lϱ����M?sZ�����A���� �7�Tg"Y�8
<��IZ|����hX!�G&�?��_�X���-�b Z@�[��ùd�X!
�C�\�2�i������R��A�3P�V��F�g*�B���X�ٙx��e��ZG�O��iה^B�;Mk��XW��xj��sB�5éx�<�^�Y�DЃS���ޚ���q�����	�%�����M��_�k?���0�j���XE�`>:ql��x ��t�������Ow����)SQ�^(��� V���q��u���������Y�JM�8*�$l�Xh���<�u�������rb�_]�Î4PϲF]_jl�^��+��c>,Hnd���}9X��d�x�Ƚ'��b�Q�e���z1�B���.Gn%!�3^k6�%]>nw��X�qJ�,���W�у#ϚL�/`��ˬ6�����w�Rǌ3�iƣel���lK.��!����v��b0}_f���O���co�b��y�x�4�2�c�^��:����ق��%&�km�Vj)so�!	;>aj�)�E������g,�m���v!���wS���^墤�����H���[�������!��C��z�G�S݋��
Ŕ�[) �y���br'��L_���>C��ѻ8\���M�~gE�K��{�|i��v����`��`Z���l�#�O9��kp9c��tc��<ʡf�a�(�r�.1K��Z$@��N�������l�����$���P{�1�nn�\��"H��ɴ�$�V��h��(Lvݝ� N����&�TG;�`��
L����n�yBjv�V"���a+jk�{E�B)�V 6���Q�v%��&R՘͂�/h���\�:=��N۪�i\�@�s۵���Z��\�JX���cK�g�1���67GM�n3A�7��*r@Tk��ܱT�����W�(��{�6��Q}U'�X�;��]��+ǘ]�׷�w��
E's�	e69=�Xnc�1�jڞ����ſ��)�o�@��r$It|tc�n��a�H�3H�Fw�C�5�� ��:r�Bς ��\�8���I^�m��Y'����ȼҝ@�Y�ٺ�#�l��MU�O�<澃�
�	d/�En.�1#�QlK��M��|]gq��?��e}���n�x�
�����j���̕���Y��������S`�,wj�M8���<a�;��i�}�}�Ŏ:��	J��k��7t��B9���4L���F��z{�p.�l������"M�'4oPA,�LT���\Ӳ+���!���@5�^B �����4>�%H��Fk�a9 �@۰�?����xp��q��^�V6�'�M-sO>ܸ�yܵ [m��٦4;�����jrί�R���/�r-ˣ�1��q;+�@�!�V��7���:Õn5��2�a<˙�$x�%�9KJ��pJvT_P��Y�U09ŧ�n�2��-�toK�M�e�Ź�U�yd���zh7~ܩ%����7�X�u��s��NU��`�b�Z���iRq��taZN�F�MI��'�;�U���x��0�m�T�L�P������;x�~�
�r{By�Re$��������a��N;�d���~��Z�O�m���#��Z �T-*W�v�	�^��
S��s��0"x4 kP��Z�LF�n�k��d�c���V .�E�[�9���^�^{S�8Fb&2Ef�z7�kކ|�!%s�V���=b�<��U�7栂#�V�������� ��5�u.v�_��	ʹ��,�O#�toMK�/���ƃ����AO���Ȝ��®3]^���u]}e�7Rc[���c�R�r�vR�(�����q���0:c(50x�&(�z���Xι�qJ�������ٍ~;h�ҿӱ�mJ��zVU㖰��
3ި�����	��
��?-�I�t�&��� ���b3j�w�cA^i�)����ZK��~f��������9�.��؀�T����")�H������U<�_������ev�,���q�^`�ib
��bLL>��"zwZ�������01[��ە������`�#���I�Om����~7>��H�{99t����9�&
��9�?�D-R��O�%q�,c*�߱	�g�����V*�4��]�y�J�yR(����Z�o�\�� JG��x</�1|!E��vh
�#9@���� 8��R��t+�	��0�p+��o%s�� ��x
Kv���ޖ{RA�B�0�f>�I%E*�ބ�0� kE%-Ż0�c��2X9XlxVHYEB    fa00     5d0�8��@AN�����;ȭ�*��%d�g��e/4DŦ�$�Ǻ�E�@��⏗,{�76�B�3��e���w�A�q�EY�e5�ەǛ9��U�D���&YA��
��J�|[�m�ؘC�E���{�J�4�j���C1.Q�[��\m{��L�C�1�ϯfV�ߍ��M�K�w�(����ﴙm��̰i�bĺ ��9��ǒ�!��"�s��c?���"����P�S��X�R�$�ΉXn[g��pKٶ��IϪV˞�ߕ�Jv��l֐��, �;�r�]��X�oR"��x�K���Z��}!�Dt�Wzh�FJ�H�n��eկ#��nC'��C��0MUّ�����������EOA���_�c?�[����P#���%(g�L��Ε�1=YQ�<�"c���2�+HVx��&SA|���a�0T�5�k�ӟ�Q����'@�2����0r={ɓ�3F�II3m"�jY�B`�D����D�@}\�u�tΔ,g���z���g�*+�J(0t]���Q�r���/�snIʚqǦƛ�8/��Cb�����zp��T�u��b�U�6`�$�eٯ�r�pr �ؾk�^#��H����Es[ >�.'��;��.D�}8��^�HXu�O�f�6�#
N�p"�!�w�f?�k�pul�7X�MN7�Z����D�F}x!�V=-hӋ^�P�'Y��e�E��+�sC#�/�j��ZZp�8*Q��4E;.D���EY��k���cf�x~�5T�aA�[]��R��"o�����dI�)��\jP�-��	�{�U�����	e:?���G㵴���g�������?\�gi.�n6�;��Y
e�w�a�[j"Qy��vo��'�m����&��Q��z����':P��W��O7�!�,)�G� �|*�<�����mmpg	Zz<�Wz��^�/T�Mc���|G+��z��le/���R�ߜJ�*Oԅ&W�(������[���)xO�E��ꅛOu@�:�w���-0R���X%Z��<��?��y�S�g��9����-����#|�(l2�H�#R}ҁlD��)�K�����> ��L�2�&𮕊](а�[���o��in��,�Ü"p ^�Bt��3F������(x��]��<�U�,d�Շ��d���Q���87,��qeQ'S�h����V�E0A�O�q�\Ua��L>��]٪u���E/�l8z�Ƨ4���Z@x ڻ���b!����wFR+$��+�S�O�9��?J))����m�c*(����}�
[�`I��{aSiˢd��H0@2������8դ��?�4�C̹b�����b�x:^Y�j�x�(�i�TR�}5n#T�a(�]0����I��,Ԛg4˒j "Q��b�鶿db\:Qpc�]s��tN�Y�<����M-=n�U�fv����2+��0u�.���bKN���
�lP���A�sN[��XlxVHYEB    fa00     640l����zkG���T
�I�&!f&���%��X�/g�)"Ύq��zcsS�R;�΢ ?-8]z��o�~P��P��e�����8�� �w{�ѾW��7�����Ɲ?�6����p\��VZ�S-��7�j�.C,�L�:��'q��Xe����+w�N:@|u��|�������t�'T�VT�M��T�;�
�3Qa(�����:_fGx��Y��Y�@C�[��:=���Ԑg�#͹�!��*3%E�uf!���Z-�K�+�aJO��ZI9E�y�[7�;��T�����1��ub��Ý��'"��y�a'��<���m�C�L���ʇ��r�
�u��O�2��~�
���ۺLv`G�1�gh�F�z�e����Y�F4W�ҷ���]�k�%P�m�K��vM�!_�=s�	P�XX��Y���"�h���y�{T�30�!R�nOb�v'j�?�V�^�[��>�|��2���k�g�Yx���Iv}��].���n<	l20z�B�K��]z�	d��9��)�B��@������DG�hR;> ������g�����U4j��[�9]���
5�F��Z-N��ڔ���u�FƏ�n�����m(V�_	�����q�[c�S�3����P犆ؘʔ���Qp�!��J��ύ%��b �FJo4�%�3�7 :�~����7�1g����ne�kݏ����?�z%�(��V�MM*�P�y��ы�`i��ef��*�v�:\��{��Q�S���}O�v|�m�ג��_�Bj��Ak[&L�I��\l�I ���� 7T����J�L�w&!�̚��`������}���fX7W��rQF����.�Hk��5b���K�(�,!�KM$" ��Ue�y ��W���}����c7h3���k�
?��̌�+�cO������RR"~u��,α�#����~�Z�R5�"�D���N��`�U�N��mB��~ʑ3�,�����X�*��k)G~�����3i�{!�D`�dn�0U��I��ũ�V��F���V]ʛY֧d�!+.aCsW�f���>	�]��I��me7�)�6��i�TZs�
�{�����Ș?x|��:SS&#u�e� C�����1pD��o�9%]]���W�©��%x��\�� w��C9�(mD'.����6y�'�A����i/N�6>�kE�SZB����jA�o�J�<��'+:�n�ۂ@˨׷ۇ� ;��c-�a�3�hŷ�����ӆ�Q�~�]�G[W�-6@U�!��ϖ���n���h���6IZ4X�4^wHsˤ��h���UhZŮ
Ͱ��-��c�X��g���R�s��z*[~��t9���s��ް�-2x�Ӧ%���Q<�
�\�X�`�$VO�~㪽�E�_P��~��.�����EM�Y���� :1F1o�O��sfd2����I�/o�y�����&+V睌3!C�t�k�m�ƅk!35�aDOG�?�pO`�y�*�ȱ���i^���zI��p�;̨�i)�,{�����ث���SK=g�q��r*7!#.��1٨,A~��[oˏS�����Ah�XlxVHYEB    fa00     5c0K��p#���u��Q�T&�P���﫫I�vLaW��ŝ}ѵe������2��UE��8Y*<��H9�����+� %~Z�ť�v�S��u ���w��8C�I���H�x���|/�`��~?�4ѱG�q�B\Շ��oT�#!kX�k=�6����ܮ2�T��ƞ�}Q��Z^���,L��ߛ�ٵe *9�sj��7Wё8��''� �=;�SI�n幀Q�8����ڱ��ˀ�Wu5]�}���e1��QO>r�5~S�����1�$�`&��:}�aϺ��!0�lJb�"ج�B�7��?Pߣ�z�z� ����_��g朡i�A�8�Ǐ<J��7�����&�6�Χ�%-`�!&��a�&c��Q%ن�c��ԏ�E�Oc#��jI ����0�Hrݑ����
y�^�*GƙE83����0D����@:r�K�� DUG�����d��|�	��(�9�՞��+J/0�6���E)u
ދ���.@�|��L�y��H!YB��\�j�z�OX4���:�.TO�T)>�Ɨ�Y��N6��tX�ϩ�R]�Hh^y5�P9i�X�r#��p�������7�(�4zu-t"s�c�懀a�����x���fЁ�u���uš�	��� �Ի��m1����N�ՋÓ��T'�.d];1��@s��.�w�{�F�Y�b����J�0z"ҒF�Q1'^d~��ϹKI��/����r(1�~�{��Д��!������ڪx+Z	1TYf�����9�ZS��\�s���E�MؑD���%�@k�.�U��	�u�)C�"}�)���z��o!ҩcb�4��z<;�Q����]�}�IQT�Rr�O���ɣ7�B�����蘆2,���XOf������"+�s�4(�TMb�ҡ�΂{��dJ���^9�����8����w*��}m��E�;ԺO!�x�*R��-4�r-�c����,r �3���N�`U�iױiT�F�������唡�Qt�\4˔�[�㍵��:<�=��Uu�����d5=��P�K�Lbݗ���'����Nһu*��_&���GWe�%*!W��J�"mO:;�'�ԼوL�2�2�" �̻��F�%�i��z����A�{�z��Ab�QT�d�b�ܸ�~�eG~��$��
c�ь.�p�w�&�7�KF�?��/H!�'�5���> n����Gz��.�w�n��>��֌�,Y�!��h
������Kgo�����ftb\�	���U����u��6��(~TV.���aK��pԟ���J��M�
O��E�v�Ue,����u���� P6W��P�ߕ2�v��.&�.7�.�C6A�%�H1�}��>��sf/�����1�7m�����-�5�`9!��N�T0��V�a��\���Ѳ�����oq�#"OxɊM�Q��	 I����]����Q���XlxVHYEB    d347     a90�3'0��X�So��6f�����x�S�NC�bj9���@���5��H�(�����,���O��2T�-�z�����B�')N�#��ޮf��\$��e�^�>�gEv�X�%�t���>��ݎg���p�A��W�W�g_e �"`��������!Q���ߊ���z|g�·���H �)�<�>Ze����z�L�>E��d��HO�V�5���� �g���8!)��(8��*\{	��`X���;�I7���;e6Ӊ��$�������2X���ä��8��a+���kI�src	��� ���+�ʇ"o��"l7���\��U,F�OR�ސ��p���}�C@ns�G�7S�!r����i��1��?"�#�x�΀��^N!��0�����D�ҙ��@Km�ʖ��T�ڱQ�}�mb���}+��w�pt�:C%i$W�-����InjЏ�O��>pY������	i�D��s��h|�`�]��Oz f3	�^g�}����"��21�6�=]A�0a�}3;?��A�Y�&�HJ1���M/82�������Vgt�0 D��dl�� ������&-h:�؊c���.[����d�r�`��6�3��|�����)��'����]y�a<{�wmZ���P��� 6*/W7��]s��;.����#�B���Ů��z�ݒ�>e����G�O�{[���� |�����)yN��@���+�� ]2;��EJ.�	�k��
#��T�^(悉A}l~5"�����Q���{�4�E���$w�f���0����|�Yv[�%� �ed��E�|5M�{w�Nx+Hm_��z�~�IqH�Y�pAŰd6�2D�\&��H5��p� l��2�;�S�eY��t�������b�g����{�
��X��Δ�Nm�u��\B��z���8^��l�3,ݣRB
~ &��{�̝~R'Z,�.��T�w'$�"
�v��XҨ9y��߻�+ <��k��f�����_�(zi�����?��q=f�����H���y>L��	&�pt*������G(��P���6+�3����ɣ�át���5T�1b|cJ��������X�!4S+�- ��T_P����ɟ��W�hI��Իײ����1���}��!�j	J)UJ��xg����7�{��@n
k��ЃlU�{N�PAaQ�;�¥�@y�O����P�X����$��8�*����{׷��9_�fF�V
�o�c��%ɀ_4*D��Ő��W��7[�}������V�{j��,���w�k~�#6n������2w+�^��B#�}�*�_C:(	�`�_��o�D�2ţr���c�N�����3 �S5L��Nf
�"Wޛ����Z��b�z����f!4	2e�^�X	�!��N;U}���j�0[��dzA�&}}��;�n��~��L���f����D�ɜC8�S"Ϝ����
]���P�mr�\k�H�
����)8w�h@i�"�T#E�A��׀���n˃��U��ϰe�wcM�cV��f��x�*�PS�m��W4���6�����
�q�*6��q��a�U!���Ǻ/��f���}��HȪ�+52B����eӓ�烏(?�J�
-������َYW20��5y	��1����g�����h;|�6���S���.�ı2��_6y�����g)���>�̘�]��Jy��Iہf"�o_�t�bS>�ǆ��o;
��̖������D�P1K���c�P��:��\.[��)o�B���s����(��5Id'RWR������>�ZZP(��܁��4B^�ʝ�q.)���c,��ފ�@<J}���v��YRl��f%��2S��WF�2l�=v7�́�E�i'�E�p��b��ɡ������@_��R�i@�$�*P�b4��]~�PL;?��OG���
o�/��4E5���Lg��U�A����Y�mق`m���tj����\��Jx�[������Řl��d72�4�J�T'�s�??��Q�o�'ԊX�hQWN>���
'�UQMXA�i\�t+��=�c�����q��5.*)#��;G�H��Jm�j�H��ge���
���/=e��:q��U�	>����md�YGR1W��L�L8�I�'=J5=�~8~��lo��өe?��[T������?-�P�� B�Z3�M��d-Cs<轆k��#P�H�1߳t%�9<���%�ֵ��pM�C�(��Y�rϒ���#'_���OB-^���ߵc���Au��x�D��{�l6���b���\~P*W���H��ՕSj�܃�o�I�$�h�S	��ǟ�UC�m���Y��
�In���	
(��dq�ߏN��z�{,��'����=AR�
����PZz��К,c͵�]�]��Vw��u��x�đf��y��$��&�UT&§����jÈ��ZBO2�kڕU8N���夵�6I��x�e� Y�\�x�ϗ��ɱ�>b����D��ٺdZ��=�?��06.c��HƩ�������{��A<WЖ�J(�3�<�/~#ɍPl�'�5 ���D?t�Iv��h. �,O:�[Zb�!��p*��*>A:,jp�~ϯ�w8��m��x�� �V5�����1`(�|ޏ4!8lg�