XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_?��p�n�n*���>uZ�AB�Q��v�ƅ��y��Z�v�ݨl� �p��op4Ҡ�ˀ��z��}��=ڎ���;�d����g�L����Xh5$Qe����i�ǃ��.�b���y����+�sf�/�����w\�����f�f�v�uX��[D.:����~��U��q��S�vG#���,&�ero�wo��X8|c��<>|��Q����F�H�0�����$����$n������x6xg�o*k�Ja�tu�x��2��U�_ٶ���g���9���|[�&���ĀU7�̩fHv�nkɾ.�vڧw,Lڷ�Y>��'���[�\�,���h�H��� �rO����E��]lོ�"oxb���9ӌ��,\Y�x����=�%��R���M���U^�ݗ�_�[U���M�"�^��0�C}8������Wn��/?� 3�cZ0�\H�ۘwz��&���y	�:E׈A�.�f2�\��-@�7�0��q�ZQ�,@�?cu�I�=#y�ipHfR���W�fL>��o�T�è��$�:֠����ړ5	��fU���Ih_��:��E7�&8ey���}X����:�e��B�P��
y#n�Ie��}@&�y���h�̋Zp���Cx��=*8�Fr��!3p� [L��*������1�7yF�j��,�r�uP-��Um��}�% ͆�5
���~����}�A6-NV�F@kJoSP���j��Lb����uk����C���'=$�pc}`�D�`8XlxVHYEB    9efe    1be0#�y��m`��A@��@�G�T���W��Fӄ�2ӭd���W_��2�fIq|$�F,EE,ܭ�cgn2��?���6A�=*�7���d����O]�.|���x��Բ�z u��U�S�A�J
�*��R#���V i)��9��{W���K4���p%�99&`��git��Xm���x��{!
�h"}J"� ��r��˺������nC��YX2�PC~��6��\�]Y�
�Ì��7G�T>g�о��g$��>{PӔk��#����\�.4���pr3�� X�+e�s��!�{?ɧ'�c�x�^�A084�l��/��[dY<(:p�,s9`�$�|?N���2��K�M��F&<�	\��($�.C��
����b�n��϶h8�a3�i\�u��r< ����8/pr�7$�-ό����Dl�����1�7#�Itz(3@�x�#$�5�
��p��!쑘r�ڿ��c���_��NC�i�,�	,�Ur^��q��'��!�
ԨUnE��^!�W����	"'&k۲�#i1�-ŷa�����y�	\�C��CeS�����"[��t���<�ʷ�K��Fq�j�4�dv�S�~_iR	�P�W��b>9;�;<-Tћ�vy�l+�I�8� cŴ��D�P?�I0�8Z�g��z�i�ޭ!�E̢�22����*�k�&KA9�|S��\U��V������Kz��&�
���lhB��|�q�$��4"=�@� bлJ��7]�v�)������{M��;?xO�ێ�B$�@��t�һ5��D��� &��c���8Z]�h ��&0�xPK�fH�X�Rw68�Rgq�{�G��LTD��;у���:*s�q�:�@m֞����!~~��8�2C	[���vn���G{�ڷ�Q�+k���=�1��=�b��*hI#�$�B���D����c��_�3��8���r���T9�}9l4+Bo���ը�,�B 0� �1��X'���ds&�BpF]�7v6p�Y�t�"[�he$2:�&�i������g�L�lF7��[��ɐ	�L\[�&�#/|>�
��,Y���`lX<}���!(!ɨ��_:Iؐ7-F�h�;�V�8��	�1c��E�Xg�N�jY�*U<~u�oFlr��2p.D߬���DI�����t��h�JNF�!D��'`��;�ҾA|y��
зi>}�SZD#���>�^� T^_[rZ�qP�9wE��Z�؛�&�u�TV�QIYO��߂�I��/����e��3��U���iz9������J8)�]������ږ.�i��l�ze����	"�j~l� �q���ZU�p�jv�} 0M�R#M`N}~]�Ѻ�dC^p�\�"H�L�H_�� ����v���
�n�C�b���_|�mh��ٯ߆�s���h�#v-�	5v�9��W�	~7�I��ч����Q�ɠJi�j�A�~�f;����z�Q�bS���Mj}-ϰ��9�S�T�|��R��4n�;���hrT�66$������P���3�ߟ��Ĉ�G��m���%AԣWκ�K;��#R����^M�)���L��#g7%��3W��E(����Z�5 ��ݒr�u���_>�/�`n����¦�puJ!����x�`:Oꡐ����$<�HI/bzF1>�x�����j��rI~���x��Bh�!�U{��S�S,��|)��"�2�w�l=I�^!�=��౒��	���HW�l�a�2��ɺ�>İ���%.(cָ�q��H�~�F��^r
�;�`ݭv!d�n�d�}U3% ߮K��ȩ>�2��V�hcyگa��{��[�m������Yf��4�[ɭ�e��  M�D')�5�禧�ɩL
6��P
<Pc�bV ��Cr  �OU9�̢jX�ۋ�7(�T�@L׿zqV��&$��R����qg�*�jeaM��Q��M�g4��_b���_�'��X+:��h�d���b��"}�:�	ގ����O���B�a�v&i����dє7)`6���/��v2�-I�S��%g|AF��"}��Eo����?m2C��%bQ��U =Þ4�Oaw��iS���d��h���̚�>�"��VPƅk'm��Z�dbc^J����z6�T~j���Z��!u�ݹ���7��G�����J�㿁�nɷOzʻ���ec@�*�Ľ���.�O������/����[	��U}V���%�ς�ϐ|H���T��BX��w��Ӭt���,�y��K%xh���L�.�%����e؆����Ѓ[�^0Ǭ��ti(�:PO�8>�ɛi�G<vp���l8�e0��fW%g�Z1:/=AVcb��e�8c�Z��H�G[{��yeD��OI䮿������0 �}HHV���E�$HR�Z�=�5U*�+.�/@�#��k�F��BxvN�L��(��ѧ���ȫ>���d�.���9yc�X�X�߶'��6��������zF}��5�*&��X�����T�A)�)o����05�Qu\{��H�$��f���a�V2�
L~�,t�l��J��cUd���%,�Z���o�S����>|�S2�9sR�V�w6 �;z�H6��<'��Xsw*�?Q��(��(�rip>�q(3�%R�!�k����{�u���K�'>��vO�Rʣ59֗l�Y@FU��v�V��ּ��Y%���-��W����]�����Yp����j�_
ի�����I�\�iB{R��0�OҾ�}��L~��Z�B
��3�ɽ*�~�e,{�(�_�`�de��O4�~4%'�T�'���ǡ}.��Eq~�t'��M�ƣ4��/l�A?�kD1�8vm�U�j�9y�tx')xL�&�k�H���O�S�(U�w�im��h��&:S�iVy���$��Q�d�ol��i(wx����L�Ŵ$9%A�=�b�>+�e`�4{��$�P���|�>��n��v	��S״\/9����6���x�[�(��Uz�9`�d0Œ+�Q�%�� ����Y�4-G%	�<���ZÔE�hf��1��4|Xf#��~:��b����u���՚�՗���w��J�#����O��~Ps�d���ܵFgsV���5�}���ة��X�BzG<F�GY��ʖߤ~����1�G��2�U=��"NR5|�4_�c礼w��K9�%=�	[lv�w�
0����a�	��퉱��H�%d���/�s!�._�%����Z= O#z^<$�W�;�w�^����C  ��H���@>]��������������,��k����N��4(Ygh��K�+�v�&��BS)��6M���X3Qإ�j�5ı���.܃���ݴ���p�1�H�-�q
Ί�뛗����N3ggS�9��KK�5�A�6�.3s�x��F�=�8�����s�.�t#>8�ܠ�2�e���Mh|�8�!(%�m��,�������Bs��A9��2f8Gz"i��k�˭oB�-J��5���n����&�퐙�UqA��Gq�؀�B�4��@�KO�-�yos�aU�	�Z�9.x�����F
��$�~�C~���R����V��>\)���fU2ҭ���N�:��7��'��o��8[ �,�U�͹"b�%!Q�[���׊�N�Ƚ��U����'��C�kn�E�Eyl��iO\�?ջ (u���Gh��������� �,��Tr?Y�T:���.@i;Z�b%s+�_]Qml_���k#�^�����}ek�tȂ1��8�!�j�ex�QVLz+:'4u��S�FM�>��z+m9g���8K�M�',|s;�����ʥ��jl��ך`Tv�%�V�;�
�#d��οke܉b#�b[m-^�bs�,���}Z�O��l�Y���VD�Kk��ό������^��6��U1����j+�Q޴�R'�1�dk�~5��$؁����o� ��6���y{I	F��A����l ?�.Z�2�~cd���^Bi�>���q=���z��+�M���;$�-
�z(i|\��1����Ч�߅�QO���[z�k�<SM|&��x�{a��xM�H�+�xc�k@�<"���\n�o)�ɧ$q���Gټ�$��ws9��@��R�f�v�;6�YY�O�lЁ��r�&�܆�o{�	|w9�-��=��d�"�\��G6W� �@���}����W�m\_�Q�g��_�}4T���z��J����&�&���%�lgt�u/w�e_�"�f#� R�i��C�u�a���`P~t��k	��`
1�[ �EWKv~M.����wI]Ex�9�x@5�![��ޗO4�� ��;��8����[��c��]��a�L��_%��"�>I��#�Ơ*H�n��m�%��K�)����_g>�˝)�r Ϊ!��wߣ�s���y�1������O�9���m$"�T��P��,s.2Tڡ�h\��@�w=�?}
s��6�q��|���>uƁ�O�V���D�>1����6��s榘}sM{Nߐ�?vC�X)L�tNַ�>8Ĉ�}��esFQ�RXPU��nuQ�/+�5:Q��Ŷ���Ϝ~w������vAN��sp��!l���ի&o/����y�J�f�������]��r	�B]�3 �]&{~��_{R<��q�KlNQ�!�a�qS>ʏ�q漮���W����"�ж�-qY'<�_k���x7㲩��nwh�<�"&c�ўF[C�i%��X`Q��6Yޣ.d��8��|d���	5�u�Ug���g�Wzڮ���V�/�C�>M��Q@�����
�r���<�`> `	T V��C���:��X3�7����9��0��[&g�J|#Q��n��6<f��R�3=���[MT:pK��r)��%CP�q���1Z "�L���=W)�P�Nb�D���g+6D	3w(�6�ECb�+e�*�4j3�*\#/lp�Y9��B��jYQh8�������mH���B���r;��$���Q!9�]�LzpC׀��t����^��|H4�H��`!��`siג� �$y�M�;щ>����1_���d�/��,��q��i�$�f���L]\#7��S=�$�sL�WU}sB���Y�0An���f�_�抭�[H�*1�����HFU0^�.f�x҅�n�ţ4�rW�ikT)%����~�ʘ�������Q왂�3�Y�[�p�F�i��_�=D:�,J�����YK����_�v6n�>X�$��o����� �Xo��	���U�9���8{3�fE�E.lՓB��龜F=�H�_M� �V��C�yJ���
5�d���6ٛ���ߏ<G<�B嫑�1�vg;��Fv�c�A��?(I� ��<G��=s�\��]|t�ʶw��8c·$C9���+`�A������F�/���D��uO�m ��Yo��%~���v�/���_q��Z:z�ƭ�@��[�]�\�m�=
���>E(殇�.��Rh�6�-�ޑ�Ǜz�׈�!��0;9�H �@xe0E�?᪝�r�4��F\�b(�)G��b���L��@`�Iblt��Y����X� ��Q3���`��X��7�Z"�U:��K��˪2C���q*�2e�u��ݑf���D���ώ
����0�1|�NG(�Bнr莋�t ����O�.y��9��GO;�C�� �~��;��j1B��V�%y�v0T�����>c������v���D��q������a�x܇ �����L�+��[C[�'�t�&X��Հ��s�O-D��}�b��5�� � 8��dS����'�Fq�fĀ�l_~5�e�e�x���)�� ��%�X�����G1������Ox�Tk�l|�`��[Qj�G�ӗ�>�����M;M)��b���
#��^��K�Όy�0��9{�j��� 0����u�����%�c-��u?��wV"ltY1"����vB��7ӾS��N�E<��)��<�mqg�O�?=#�h�~	�;UH�����[�ɚ���tǜ3�<���;��/�kϏNK)X�W����\��!�Fp����Q�\�p�&D�K]�:�-�W����]ϴX��.7���0h(�����WQ��t�Y��	� u�8�F�~\o\�F�m������͑���	°v�~RɁ�yW��M�7K�Xz_�ʲ^�*�1:~�&I��	#�*�O<�c�jr�"�� ��tZ4�"j���xO��'��V�}e��b���6���$�^]��I��#�+3�Ho���B)����_~J�m��������0r i�[WKY�E�A�ހL���~��9�84Vֻpҵ6&tEMO9��<�V~�y��^o?���ހc�U~^%tC�6�+�T�򾮋0�-2��T�b�ȇ2�)�F�TU3��t0�Fů\ʃĲ(,��5�ϩ�μM��6L�Yg�X+�5��dQ�t h���6��<.�腖��BL{ܐZ� �b ��d1ԃ��չ�EU���\˓p��z+���o1 s\WdC�3��9�����V��&�+����t>W����mXYЮ3տ�"�G���;��0��@br���
�!��ɜ���e��ǥ�x!�s�+3w��1ϝ����L~-s/&Wf�`nɧ��%��_�ݹ�{�Mhc���-�|'ڞ.R�ok��`��NF������!A������^S��D������V�{Fe��2T��z��X�9GnM��Wl��x;{X�Vdw��FD���Օt�K�!A���UE�r�0C@p�U�I��\u���P��*����?Z��?��9��i�)�;�Z�tb��dF��
�N�:	Tt�Zh��E}����u�%�MIJ�P��X��"�]�������u�������ʫj�>2��=9�1-�z�1�:���9zr"�]��Г��P���`�0�}y��\�>V�8;�Y�����w�ҕ�^άV7��c3*}��!����	���E麷�d�t���1���o ���1�`���wԵ�i���w��`����7�B����J