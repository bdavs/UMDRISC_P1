XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\-$;��,���9Xo��M/�x�ն���e�N���|O�*�/���lY|u���6���"��Hd�o���M��g	I�����`aN�)_I����)dl��r����`<AXh���9Z��[N&t޿{��P��0����/��3rT���Ƕ����� h�x�7��� j�@�Q��2���,��^w��R�U��FΘ�̻�l�h��WyY`��h��J.DO��gѨ�mI�Г�5�4���w<#M�t{��Ad#�A���4hj@���MW����v���O(��������Q�t������ne)I��=�ۇ�JYau�̨�	�&�e����uS}4��P����s��D��Je���K%mmeʠ�2�얐 !�1[��9�|Ԃׯ�`Z�Q�ց�y�D�u��"l���M)L�a���_mG�?�639�-�4l�0g�)X��t
���OAĉ]��+){�a���HT���}I������ ��2��W4ɸ�Q��p�:7�a�[��]D�����_д ����_�m�&�ęѲ��YF��Q�u�����/
Ȳ�efH�cFMMD�>l���;a�C��)�h�{�����}6�NV�Wg�.�2��[���rh��}�[�k(t!jA +�#`�}�U �5���5lj��c�ܐ.;ip��PƠc`�J7k?���ۂo+�� �B�E�/��*�S����*̄�.�B4\X�hl�=��X\�!����-���XlxVHYEB    fa00    2d60�<�d��O����kVF�,YN\e��c����-�y>0������ �R[	��e�_H�i�n4�R�/�G�S�9����|�Ƅ�"ˊ�������wn..5�ea���X�ɪ�壟o|�ӌF[0%�;����0ڠ��]�=~���
�zq�R�u�#^����I���/l�QU72*�V����4\/�/��A��>)����s}����6Ee/ qHe�Cٹ	ğ!
����M�c[z������ĿP9�2��4���9��l],�M�4��LCܙ�=u^�θ�TH�	 ףq���>����:ְ�49f�'�x�Rb �����p]���Y��!n�� ���	�7mG��g�r`���"&�I���bÄ×�\"�6����7����1���N5;&�t�j	�eeT߼p'�������o��%��d(���J>72^[�o1�ZL�d<!���~$��[�WT�8�cyr"�*�ߑ@��*K�C�|1���!��6�km�`}��sG@y�aF��y���C��)D��KL
hh�}T4G��Ƽ(�r0��;QF����U7�rG����oE=���1�@t�w�t�e%K���z�7��3�=��?J��,0���+R��3�l��E��P��"�/-��L�$��N�-?��-�a�qN�kcF�[&����RY��*1}n�;-�5���@Hc��xA�}sAl�U�w��<j�aB�UUmM�0��H�7�7nq�\��C3ogU1��R8�#�<J`?�BX�vX�2�+�wI��uh�M�b��t��_�iެ���
��1r���G
��J�?D�kˏ�
��KM�YR��B|U�ޥ�Ƌ����m; vv�S��O� ���"��	Z�N'���B>����d�)L�N�U�eC����f 1i2<�Pr��#���V��]w-";9W�:�D����m�<�ɡ��;�غ`�����F�+<��h��+��z��;-UN��o�E��p��	 ��ry�ce��|¼�:<2�2OX[�� �IX��u�V�k�0/w�����j*o$AɄ
v�Ax�=�N��� `�x��>�L� ���'_gm�H���*��љ��DwJ�B�7��%дoB3A7��yO�Qw_�o�#[�EC���v�y���:?ȱ�9�6nD�A����
�.Bi�R��c�Y�Mc��U�d.:���+y�|�VhF��y#�7�U*�+<)9} �-%�a/zw_H��$P�㹘3@��PhE}��B��:Ӌd�%���p�<O����xX�'�������<�F/z�"{���R�Mn�A�[2�o 1�Z�ѡ�z�/Th����u�k��\����B���:�b�����B�Nƽ�c�.���5OL̈�u�B�8�k
���_�+0܁Ϝj�@�+��?�V�.�{d�T T3���n�n�P둇�1JnP��|�GQX���\������&�<�U�L���Ws���cSԽ��ö�����\p �J��i�>�X��\�L+x�;9Jxp#���^�w�Us��ߊ��˨Y���3�y��=$���Y���UI��>p .�i݅�	N�0-P�e�my��]�n�
f���T�*����[���V_��+����x�� ���"�${���r( r��#���?�@bLq�x���A�X%S��Oۧ<c�GlDxX讂�.ڻ �B�>� �-C"������gS��:�W��!3�W����gK	sԤ��޻�����[�.��J}pk��y<g�Kr��U�zԿ�7t��2�'wL,�@���X�w��7nX�Kf���a.�8^����\�)�G��$��W�i%O�#=�]l�P	"d�ݛ��h0@�TL4˘���ބ��J�.V�ć��#c���;��mt@� �c��Ē;�C�2����<��n^O�{U\Xi]F��C��un,��Ǒ>��БG���9EM��v����|�ʄl!Qi*c�5�h�e�����L������5���cAoU
l��5�&j�+r�$P�0B��_��E5��O��_�U��zq�đ���H�9�4��PAł�+�����9�-���3�ǪC�h�I���	R��'j
/��K�� 桚9Q[��7���N^�6В=���ߚ NT���s[�!���yK�P�L��ć��cŊy��͛���������6 �i.!��D���0����,��j"ELwjR����!8�4���qn�	�?�,�M
���&�Qz��'v.F9��	��<��=�ϸ��6�*��{� ��j�����o��pU���i�wj��7k/�� ��r��O`���B�閲vV�X�ge.77�@w�u��/9����cB ��h����l,���q�!���X(��N���P6g]�0ւ�.�����L���F$rbrW�N��^@h�q�#aQ;��}�l�����R�`U�:͊0(b��t�����~�j�"�P�E�j�KP�;�5��FI�>B}c�fܐ��i�S(�f�l���z y��xt��)��i��+��ո�h�U䞫����B՞�ݤ�t�6§3��Y�*����[�A��e�as�m�2�D[��ĵUY����G��d�}7>ڶY�(�b�-�)3/����0ʪ)f�zr���X���I�������ry|C��^�V4���,�1�ȱ�"���q��EqA���\+���<�� ��(xb�iI�6��s�6��jv��G�!p�Q�WkD�W)��R�A	쳂���6NAݣ�'lUcP%�z��p�(5��a�F�7���/l���:�6GB�1L.�1{vV-N!�9���L�F*�nz��Z�#~8�"!0�d"�	`�K���R�;q�n��wў�&p�9����y����,˷5�2C�g�������S�g��֏0O�n'Ju(�I�X�=�ì,�"�ꥋN�� �NwL���ל����sC�K�#����-�f��y��7���fH�g�T�|�K�f�P�jH������M`��������b	�Ӥ�AמܭV�s�):�o���R�,�3W�T2�w�o�tA��v����\TN]�o��ȝ:t�r4�L7v�(z�3q[M�e��sR���X�&�)�G��Һv�s���"o�����2�a�pHw��`TD����x Z֥�d�J�7����;<& �\B��1e�Z2=�n^Igr�I)���&Mt���r��U���]$��[�Ɛ�X�u[��tz?#���A^��2�����K��1�Slj���A�z��$L�/�����&r���٬'���
�E%�R(�p��J�]�!�����]�k)�T���,	.aj�p������V��@��/����Jf���ne���q�_&�@�:�]h=Z��/�S�8�X���E�� �'Eh���(\A�*���=r6��010��Gv9�Xl�p�h�����o��}���?��nZ���ץP���!P�޶�v��c�"B�n�����#��H�7���z��{�*�eq�1��ㆷ�s.��%o�
1��&��ڰ5k�K%���.v�Q����׺�2��Q� K�*4^e�2��(����)
0��®��,t�j�P��o��&8z�nR�P��
�f�p���=>�RQ[Vu� �T�0Z��V��ƒ.`���{�c�n�-M8�+�bir�O1d/��kq���o����t�������D�:��q�4bA��[���͝%�?�U���h^8E{�Q�l�o�h���N���G�^��i��@Ҟ�~m�B�.sc�o[`�����Ri\�Z >!�җS�2�E�9��<���T����0I����w!�{ںh~����.�S�����ɻG�����c�i�� �z�4R@�Z!�Q�u�:��r?'�9���	�4O������	��V0��#� �	��QM~`����"_CO�\�jX��~��t+4�r}�r��]O￉�M�KY�t��B�?rH9K�z@�3#f6q���ǔ	�;_���o�1�lq�������Z�<[W=�g���g���}����J�����B���BX�+=[���R�Q�?�ᐿ�wE�#I�@�2�y#��B�x8
���t�xy�9LM���Y��n��T����Z,�Ux�S"6O��SJ\�3��(��|��澡U�)2��� y�9�&�Z�h��D��x��͞'�Ң�(����,~�F;��86�[�xw[ǅ���?�/pL�l��q����+{fA�i��4�y�m1�����idA���a_�}��������y-Rxd�h��Pk��>�uo�z�	�]F�z�mf����b^'�x�<�Q��U�����k{��e�z�$q�f S�3���+��(^]�LϻD��[����l�HO�^B�o6/~K80�ǫ?�^��[�&W�G���*;��7�Cr�����ӎ����n�I���k����8	�]��ىs��T��c��AD"Y'E@;��*������dO�����|>�T�)�"�g�(�X�Y�a�@�e�w��3p\yة�\Ԗ��f>|��z������K1��5�z=���0�I�t���5F��0�Zy��]?NBn����-rv��l���Bo���4 };��V�͖�����뷉��}�i�#��4YB~�mI�
.5�g�J�`A~C����LL�EF/��\��Y��n��hMr�O-�kf�����Xc��ڮt�|l��6�Z��,�ǎJ���\	!iV�
o����̊��T��l���|�	�����9�&���gϼ�]ӛ�"Wn��?T����q,�����+�%�M������J/�5��7�Qugt'�Q�
�^������>�{�p'9ſ�U����v�筤p���B)���}1�KE�><��8Ҡ�,��"�4��L����*"D��C "ە&I-�e��ٶ3^�,y��Y3�\��\�[�i��Mj�ɉl���eP4��{��%윿��l�����F~v�����wS>�M�4v¸
�����#��*� $߾��aʩ���� zq���[��!�n��1��w���m }a�'��U��P�N��#uV�{8�)QIIb��YJ�G�5�<�������Y�$[Q���0��p�{;�r[���4c��'/*���V4���s�Z��<�)�!�g%nk4E�C��Q��nH�dn�
��mm!Hܲ�}>
�V���U�Z�_�+����VQ�~�E��K7]��6;��v�;mѿw �+�H�__gc�4b cvZ�	���+�u��kR��$EK3r9R�g,�O����FlM^�Z�F��o�qcQ~�.�%��zH/p�jY�������}j1ǓW���/����ϹD�N2��i1D#��As[��qe"OL2�>����-:NϺG���Px�:����f��>���\�sֆ���=�Ā�~g�#4HXFՐi��V�"⇭@3afa�Z�Z<��B�aS|��E��p�ɥ��S*����W�>���T��S�����U@����0��3��4��t�/�������Fp�+�!
��h��������M4��M�$�6��Xd]!X��zKK���PP�T��0嫁�U6�n,��v�j���D��r$@ow��>� �~����7����;��5�R�k�{�C��99EӍ$}�����P�c���[-5����q�!l��&>n����}�'�s凞 z�^��ls�����&�J2�>n(MEi�́U�z��y��=V�[�l��`{���J�ʬ��*>�!��GdW�90^��1C.eߖ���坶���OJ�E��ڰ�D��ń*8�#gŬRf�
4^�Nc櫒z,�r�p7kP��MFzz��K-�5�pi� R��I`c��Q����"7�LVd�t������Z�¬զ`/V�C�?orq4}�?XG�x����i��`�IhA�'ͣ!�BݩYy�x8�R�M���Ie�[Q�}�k�!�Y1��y��3Zً������!}��h[���:;��Q�8��H4��wC��$�;l��Q;Vq�.[���^��,[(	D�:�b"���%aE=-�;�<�(Z9�i������u���'	�$�H����� �h 8$佉�@P�S��KE�,�p.�=��a<�י�=Jߜ�n�	��Zc6��3�gC�+cR	���tU�&�{�k���r�w����g;/~Ěj	�h�S�����͔�E���pC}�A���:/���u?��l�_FE���I�o<���cg5s=�K�Ud2!��럂�Tqf�� ����;G��� �k��1�?̈�]6�>@0�N�Z#ls��٪E�)=�A)�Ҷ�y�Q����f{#�Ѿ�c���\M�˞EQ嗌,6:�a����N�!�������p';9��,	w������6��B���t����r����̄����X ��}��D+Keb.e�g�l�c�%7����ҲP9W�`����HX��C�D�.����ae�<6-�y�;m��6�[s�D�G�҉ 4��~v��� ������	9p�������Ҕ4J�)ŀ8��W�@����
��EP�وM?5������rA��A�(���{7w`2@#�'*�u�GϞ2z��Tc�V�1$}!������ñ^���h�/��7�q�vP�Jg��9fAe��$6�H243����
蜼��W)����E�j�x&�&�E�o{N��Xmk��"�ki~�_dq��s�������&Vﺺ��N�2�s���q�UO������N�ɺ,�pP[G�Z���.Ql��r=	���m��S�)�tiz�'g�X#Vb�d������#�	�/{��]*�O�
Š�J"<P֘�1��%��y �r��Yh�ޖ�UУŔ�4=�������k���?$J| M��{@5���\S&8o���:2+=�ڱ�H��мS�Y�#��\�{XM"��>s��j:4q�4��L}�+�U�]5��+��?�K�
*�]_6��mS����r�aGx~K�LuyN�!�����O�Qi���tC3O���-��0�'mr,���p?B8I�-	�,��cQ��@��G�����
�Vv4����U�!�0�➟Q�W̙7�u��̢�_��(��1�+��V*xً���_j〈@'�:)��jvf��$M�WǑ3�+j횘�K��\�8@��nʋ�6
��aN������s�m�@�&��D�J"d7�dҫt��$�W��9�Q��1��hj���%&���eM�{Ɇ'L��-'H��!�e�!Z��ɒ����p�mU-щ�QY��j'��i_K���M��U)�q��ah��	�����F����B�90�P#��L�^�$�2ۦ� �9��uVa6MZ7(�g�������'�4R�j�]���Ĳr���?M�wi�):�� �K��̽�63��^�ͽ�2�c��5G� "R�[�v68��)t�;d�!���W�̧A tڼ����T��A!�����cԐ�Ï+B_�=����m�=k��m �� i��Cg"�h�8!����"柍O��8�IJ-.�fS=VPis�%��2*l/LVfp^�C4�襟������:�t��0���~�R!LiyB��Z>	�k��z�� 7��5����R��@�49~&�����.����������,}c�l&z���"����APԷ�E��:��{���$�FA�Fm�[�.��DX�c�rυi�7M&ʀ&�v� �郖a�p����W��˺}�W����}�����蛣pjN
�݋u��$�����+���WFY3%YR'��Pu��M� �)�y�=�^��jrU�`�R�o6*3*���AQϴ������i� r)�A�/���n)_z&~��G/��"q"Q�=E��0!�]�,	�ly|�2�dg�[�ࣇU̩0��rv^S{,�W�X&E�L��=0h���d����X�Y�gK��I�Mp!�:t�,��SHg��ݡv���n8�"�޸+�/�_�S�	r��S^�p���!����4�R��֌��J+	��#����ϻ�]���%]����U�p��5�xV��h#\�D��fV&�UZA���B���۵�q~cN���wm�]ӀrD���
&~�e�O�3�
;nYs��	����(|t����;�!;8��PUD�듽�Qaт!�ϵ�	��y�����8c�:R�N3V�YT�"e%��
�x�?.��/���w�L�d�d����1���Q��=k�ٔӈ03�Y����7)=�:���%J��k|��-LPl��e�S�Q��ī�6<m<~������	�Ԃ�d��z��k�zUӇu�����q�O�{�o8������á�q�	�0%�IR�&q0*V�p?6v����4oWN�T��*kZܝ@n:����7���i�|�Oܚk�2"��5�ZF`d��������ݏ�WқL�$��)��hcX�杗�"��-��]�<b��� ���b��������C&^Yh֧X��T[_�=���*�a8;��r��g����VL W�� ���?l��/00�m{w �ހdJh@�r�6+b=��#�4��$�L����$�K��	Ê����/�u�HY.eB�f���Y��~��&�/��5Sqa��?Y4����8�y�<�S�<P~�@�V��,���GK��
P�#�rt�撅C����!�N\q>	Wo�/��cNk?SƗ*:!���R��zB��J6�B܆v���F��ҕj��px�m����A i��R�֚�W}�n���j�Iq�I�R�0m=��Z�����3�-�������S=N�����45Q}�{@����>�*�,$��cr�v����u��3�A�!y���V�#8�B��i��H�/i�-]�~��$�5�{���rQE����Զ"��P҄,�'��L�9���k�N��~�1�D�U����������KI�V<w�����p�T�T�3fM�G�+�JE5Lj��(UI���zI����=��w��Պ6v�7a�,_��
��T-D��3�-��R�s]��k!W�ǔ�WO��E�膇1{��8��|��0ƥ
!���1��@w���m!��0@�+�dR��w|*�h7�x�f������e��̒l?�M<!7/������p=�Pʅ#0׮��:�1�-6+��'����Z�k��v����VL2&�#�{��m��ɓ��㌠����Mc9��x6C�0��iXj�1�&,wZl;����=\Ǹ�ؓok�5�O5)�pW�ׄ��Po=����ڼ�����UԵ+���~�}�2Ǿ���$
�U�?��t�XAZ�ͅ!�a�\����h7�;�IH��-��p�bMw���C������uv��)U�/3�=�]{NU/R}�hA�� <�v��][ߝ�<��ŝ$��aN�I��Њ����L�_�/<�BM-�%x�C*�lS�_�8e�3����^ݍR������"��~.��#h���A<�P�u
���z�g�	/�B:$��7�B<�XvU9F`�����}�ͷ�nx��#t8�:���Z��6^��e�R:Ch�E�DAq�6�D�r1�ڄ�ߦ8�4*�;��H
����-۸�8�,��#��RZ��c8-C,E-Ѫ_j��4�TR��*�!�XCyZ�71152�m�8�F�iR�-�	�s�J�2�%m��׈�����?�y�Z'��8c��}rdt�rlE�m��6f��8�_�⨗
�9�8�V�̦H}����aS���v]a�e\��v�RzM�� H>cg5�{��甜��}ev6M&H3�E��܎ϏxY��V/x	��U
m�#�枍`�T��rןctQ�C� ������O8x7�Cs��K��"��GV�}�?'�.�����vB�i��j3��٢r���:��p��rK��k��½�/�z��Ջ~I|G�����=�>�҆�GƯ*'�5u �>���@�贴a�!~�{��fJFߚ�h?�/n�{.m�]��n�f`���%u�� ƠZ�m�A�[=��{ċ
��ܩu�m���氀B:�,wB.�;V�DK�����#Z᯦��6(��4�i��G�V�b��*�����1�:Zsܽ���d����ΎN�v��������~`���{L�����5��G�gҪ�LKݵ��v��ן� 
��$���e�[2�%�K�NJ&�.Y�o9i���c-{u�iW��ļ�գ?R
��9s(dF]�[+:�ܦ�޺ܫ���ҰԜ�m�Q{��Uї��u"��u4\yg�a��:��R��{�i�N��b�L+��ȉ;�Ѽ��͟�tj�EE<����oqeq�7��k���zt7�(��,Oq����3y����"�+k�m�}C$7�M�fT�ز��n-K�ƦS�	�a� ��@���0E$I����!�'ҧW��bG�֝2���7�1��؛�(I�A���p��X._Lh�X?-���q��H�FS�����a[�xdR�`)�z�F;���v��_�FF����f*�E����h�o[t�Ϛ��CU�]��2����β(�rW�9����l^qX���Xױ9�����Q���"!Oǜ��K��U��q7�˕����V�|����.1�?T��ᆞ�9����t������7�u�N�I2�h
G��,܊���G�.7y�*�N� BU��'ɥ�����F�5]��!��Q�V��
���LHJ�Vf��Up�����u^���M�K��L�u�+��F��`��Q\㨡�7�R����%���:'GH���]$lm�*߭k6�M@�p��$Bi؃(AI�{�ˑ�=�Ҫ�9+�o�-�!#`�����K>���/�����4��X�Ǝ+�H1|�j%(��у�X�!.��1"�����-���|�!��@5d��J�s��1�a%��%�u���Nz2'�8S͎��&� ^�%,�
q��mWuc�M ��������#�ٓ��G
�̏O��ROjN�׫�C�	˵�d��_]7}�4\��.�I0��V�P�Ɨz����CY�IY^��Y����k�r֥�y�?�"�{��l/�8�?�/�]NԦ.��l�B�ܧ;X����Eq2I�Tq���C+���n��+VqP��tq��B��选)������.FQ4V1vn��R�y��֕��C0���+3��e�S�>���A,
$U{�������gD�窒V�恾hb)�t�'���5�?]R}0)s�s5��þ�G��"�ʴ�C��2���&�:�(M�V�c�1V��x��x]�V�v���|p��@�H�`?,HE�K�������Q=�H��'��4/A-������ҦWdGZżガ*$�H�n� �x�$ֳ��=���ǧ"���X;c����4����P�/S��v*9!�ܽ�*���XlxVHYEB    5914     f20k��!s�L�����Vw�5-h�X�򷡅���Ŵ�{������b㼈������Ⱂ�al������E96�c+;IGr�GJ�qY��e�f!��}� ��Q��z�R��H!l�虎�'j/O`)��T^G����ē�E�4}�Ѥ�ȐL��4�$j�|��8fcŚ�������+zw���HUOfL�;���S#�����ݱ�l/X�Q5���{�W��n*�v���ٰ\֓@�b�\�����j��K��[h '�[���{��JTE6Ս�p8j�@��-"��U�־�(�/6��GH�Ĉ�;�Ñ4�%�I2I{��L^0&�o�班�w�r�8������&[ 1|� ���X{��afz	���$e?l\�RD�f��%�1J��a"�1�7=Jѣ�����}�+�׊�8H����'�o���0vhT�pP7�5b��L����=��)Co2R��!�ǔ'd�)����P'~I��);ږ����;ĺ��/h^��).!l������ǹ~���}�~��'�5�b*^�D&���E�)o�1t7�E;���.���`��	��s����l���5` )4�����Üv�
钲q�	-ɥ;�����AX�쀪k�(�A#���W���:l�2��{��P���'�/���n� � õ��!$F|� ���95��Uk^�`�<����1�,�G�<��?�SyM%)W�"a�*o�~��\�^Ҥº}O���w��ҫX�#E���'�\��oL��u�O�뤖��5)0_����LJ�m�}+�� S�[�����ݛJ,�S*ޜ�N-^m��c��9й�4�˙�����4�8�֨�?��0�D\r�d��j;�e���\���k�Fl���T+�i�N];� ������"8�I�Ļ��>py;�]Mݜb�aԒ��ԥ�n�*4�B�R)G��$�| 4&�]xߝxm?�f
}�d��b�O>0nl���ӇLI��������ϟ�<R!��- �D�ѐ#8��?���I�?8K1��d��!i<�!$�bn���MC��z�so==m�o݈i��i��R���[1O��]���dK�����_�ז�o�g��Yy��F�̽��d���۱��I�;���1�*�Yh��@>� �U��*�c�܎�Og}�|HZ�{�6V���(�f؁J84q^��8V��"n_k]Y9�԰Vkjb�+��Sl+w0T��{}FCj��YJ���աG�����<t~B���G�S��R��	[��9�ȤP��,TRg ]=��^�n ��.h]��������Ȕ̵_�Ui� ):7�۸yWF8�L��%;�o�����gpU*$�^Ze)��"�C��y��\6���R�Ү�b�q;��$�V-���r�}Ysӄ/�z�}v�@��Z�h��a5[]�ϐ�F�����-�����6P��[��k����_[;�ԭo%��l��a�����׆e�"�Y�Ծ�q�1�@��V�$�b&އ���;�.��(Y=��>�
�����Ð= �������O�u�����N�Iҗӌ�s�9z���a���Vk��d�#~z=�}]L�ۂ�����̘W�A�H�ԡ�j���8M���"�*���l"5%�7L_�]���+��]sv|��	��&�Z=E�-5ژ�&�kzi�9VD`�,�3��׿��@�*аo�_k��	f �M�/CJ��=t*i��5`���om����)���������ʍ�C��3���gK�mF�߽T�������%�c�L�T��lxiﻚ���oP0Z�����3��8��b��������Xf
�O�``�x��Dmi�}���N��Oš�X)���Q
a����m�O��23��F��T�;˲Ű��l��	���\�4�W+�(�I��1��)�'k�Y,�����uM&®}a2�����9�R]��Α��C���rV@��J�"��d'E.
Z�0�?*;,��M��Ig␈�N
mp��2n�S������Cb`���A�/&��j�\'��DZ���C����ɮ+��2u�Ԛ��7���4�=a~ճ-�RY�"�;cW,b�1OD�����[��J���������b�f-�D����y�T��>����̜ݍ���8�'�5�]PC�/�ƐmR��.l}�5X)լ������'�+_�.lq�C�8� WN[�[���'�e%�JIuMt�F?Mw��u<<C�Υiz�M��C��t�*�L�OkI�Legnv�F-BI��Ϩ�<ѹpT��Ў��YMZ�+�g��oW���P��g���a��\��$u�@���fܨ�j��b��k!�+����I���hݑE��o����܏~$�e�����硳v�����K�Y^��ŭ2i�W�����p�h�k`��Ey�u�;	\�[�B�{�}`mX��I
b��\�W�z��#7��~�a�-���ՏrD�;/� _���� �_��ӟ�<<�tXc�*?�烗����ጤHI�|�s&�z���v���ėW�a$�Ⲗ5���d��X{g��t^k wS��'�E�`�J&���V�_��Z���Z��q}YXc�	��F�`�w��-��T6 �`z-X.��d�u��������#��E_�.�R�G|!�/WÂ6��dR��\����99o��X�������-����)�ov����{w����+�W[�
���{*�-5�rƃO�+{Lmud�I�w��fm>�A����,��aC�%�fQ<S�%0:�<�#M�xJ��-��Cx�X���+H2"e�r�����h�]�ķ���@��O�Ge�Y���Q��D��cF�.]eH7�s�=,��A����J͍�w�DX��ŏ�t3U>��x8Ъ�<yb ��Y3d~�9x�Po�,
��h|?��P1
�#�Y����ﵓi9���V��y#߹��8Ŭ8i:G�f���Ý�d��[qu�:d��2q��Y�l;\O�yg��]�y�Y�w�_�K�c#�
�{��n��@g2�;�/Y�9
�\w�f�������
�.-��;����L�����J������E0�F�+IX�r�}��JY�~��5H�nE7Y��O�}_dEv������>�&Q�hõ��t�7)�|��y�S��k`{��a������`�p"�Չ�Cٟ@s(��v��kK���ղ����������G���-$V\&���V���*���B�+B	��T���%�@�,�.�R��A��텼w��]b[�+�k�1~h��q7y��5���A�ݪb%<H��u�������x<�x�mj�:Wc���=��e֟�m�k �tӠա(ǌDj��YJ��ٴ�{��䥔��ۙ�WL���FЄ�y*�1���`���de�5;�~�������)�x�J���iK�QW�<���Y�<M\��{��Ĝ�����y]��k�!���� -��q�N�����p���I�}�\@J�oW��vRnq�������P��˿�-{�������y������	Hg��d��Q��h�)}��K��m�@?��\W�`jߙg�xd�QŞ�I;�"��b�o��{nz����u���)�՝�E���ݲC���39`_�M��8�A==�w��%�EeX{&B'�ٖE�V���,s��}gyԱF&	y¢� �l�k9E��*+y�2�h��U}�^���ƛ$_���0 ������[n9�i@���NfX�	_F���
_E�g>�4���[e��p4�_C�qJ��M�^Ծ�?����\f����