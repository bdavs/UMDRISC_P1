XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I����}s�i��)����׶� 
�%�k�np����e�<�P��q���A�+f���a��f�Y��֙�u�J�:���qa`��@��`++�����v��Ť�l��pc@bޯ,3��e����/��z����"V_F	��)�h +ML���u�=�R�s�[�
~�?&�|��G\��/������QA;<w[H�-�;t$: �F%��=[~�i8a`2��E�3�.<��jtr`���[ZI�8їw4D�p!�,05E׼g�z4�BwX�3�@:?��n-a���t���`��#r�K}��-�"��QLB�����,gČn�7�������ӌ?$|7噤�N���G$ǉ׋%]�uyV������'��S�>��Rr>ɑ�>nn�	�U�9��(>�	����g�8m4�AF��Py�f��$pDAl>-#����$�ib�=QO�[��+1:��WҝC�!�e�ڍ� kؘ�"x��[-l���4��pS��#�ʁ�,������k��@�	�c�ʨ��z�p�L�����Gr.̳<Q��7g_�^�m�cbA��q��޾]��ƻ�2�z�� Ì8~U&���҆�#�B
�۴���K�q���v6�#Oͧ�^H:�%�,��_*�U�^�oi�n�AFc!���[�6ha:ӏ��۵҅��=�`gQ0�YU�����_�����-v�k��Eo0N^w�����h�^]�I�ٱ���ϻ���Z�j�T ����
;{�Q��l�ӞȈ���>���ӽXlxVHYEB    c3e8    1d20�����������_��y��.�0�wkJ{!����C���2�T��	t��7Y:U؞%84��I߾�@��:�C�����C�t�i���U��<t�S�m`��U�4�ۭs��W�9���A�d���42�ߨm�,�궒T��26�ۄ�*�_��`��Y��J��e���7�WLg��6C춏eT!߄5�?aN�6oS�
Kx8�{�;�G>4�Zv$� �v�%�U�A��柭���f�#$���x����rq|����^Gp?�BeC�sn�=?�o��ě�T�>�}�(���/���������M*㡑\-{���>Ec�H�1#�٣�R�7��+�&UXnՋ.�%'NlSmr9dYm7AtHFG��p���{�[/�|s0��8�������`� >Z?&E3�L'ݙ��3����1o
��u\r@\JH��XRfyw{�n�v�8s]��h�/v�R���i͒K��I�i����g鈞�{*wTRi�ڲ3� �K��aY�"� �p��oޤ#̉6���s�#�(�w��G`b���"&숎�y6��$c�^�6��1���n�O|�U_ȃ)s%SxO<6�U���ek<�`�3c�˾UQR�i&j�W�=��f�V�<���u�9y�u�lr#�#��_��ﵗ9�C�^I��שR�Jlz�j(��-9��r���Ǡ�]�k�T��"3�P�����6��%�gڌ��}}�"��#G�K6�SD6 }�6a�C.���EK��3H���th[�u%OsL��&-89�ԗ��rP�AV��<$�A�F�vZc_끴��ʘߘ�)=�\0�۳h�(���Ig�R����yM���A6����l�Dy���r�jW�������ړ�4��L!P)��n�J �\}Fw ��n�&��o��ZT��� l@�'���XҠ�� ���G0��0ݖ�[���#�\3�3l��_�Ĵ����B}e�`��&֧��A������ە�y��zM���Y��\}��^c�n�*�6��� j��ǣ�e�C�c!S��������bc��jrlx�*K-�0��ʿi�f��s���P���s'�`ܿdl�'���ֵސ���i�]V����t@a�Q��1�7�\�K�R���f�L���4]:sB~����^��'��Qi�ķr�����_	�l�Ō?�ܖ�4E۴L�c,�j��o.��+~��CR����bYGn��9!$�����?#��h�@R!���zh��6����>�L��V�rRS�aP	M�����7�T����T�,hX備�1���?�K*�'����Db���L�n�-&� �J�Ɏ�&����7�2nFz���6��[ �>��U���N�W�6�=V�b)���16�%±q]�rh<��V$?�#�����zg�!���_����3�ۮ������O���'˽O^�s�qp��nSY��}!��ѵ�� ��M)v,���-@O�D7�XV�!ld��mg7?��Bp0%[�5��̀�E�p�w���*<����IN�*_�_#���k�1.�Fhkă�50�ڡ���έ�ᙜ*Jњ�����*?��MA��l�����./dF~ۘ!�#�zW�V7��%����М�;���٬Q�D��97nЁW(��k ը~�M���G���ح�]�o��^I}��n�j�f�.MV�GhK�ZM��C�]�|^�h9#�=gL֜��}
��-�AK�B���&���؞�bH�	�@�߿�|��(�$��T|Џ� �/�ݷ��=��H��)[�&ym3,���C \hw���r�U��تvD#���n�93j{Hr� UF	�	�IlHMX���h�|r�Fw{�i��6��W^�QMY�p�r�W_Z//KY��6A��8����t>	��fy�V#�$8�W*c��L�2�a���o��},��(	�ܹű|Q�z��+J2(Q�D����h�3��rr�[:��P��u�bn�?��]��|��@t�V�ݡ-XP����ʀ�q�{��s���=��)A%
m�߰&6٣FЍ���	0��F�0����Ҧ1��'X���x	����/s�ߤ�EH����D�(�b����D�)t��3�!���#����L2RV�0����0K��-3�]�[�j���Y띥����C���G���O�|"���Of`Xcq�:�ץ:�xz'3�����]���d��s�S�7{i�
c�C&��I�č�0dˉjQQ���\�<<���S[��-��u�$�B��2��}cY�x����+��0�j\� ���_����5���j�A�����n�Py�D�2b���]��=b�Dj.˳ۍ\�PF�n0�f%Q;{l!t�ㅧ����SAυf�U�e�kZ����S��hd�\��G�i�P�l��+��	��/����bޱ��+c�fX3�ȍ1~���vGk�wo����_�E~�'�ߊV	�2a]�+z��N�&l7���d1���.��͜������NR`�*�Ȫ�KG�϶��kk�[V��i *��V�M2ځ>}˺��B�:7soOlJ��g�;��FV��͘��a��r,k_N�з��B��"7�9_.�!�P�-�fc��(�k.@�H����&Kҁ=lAs�q8��`���LO2��JHC��ի�`��h ���eK���6�
3:�w������z<�LuQ��I'F�Z_1I��J�oXʼ�BW@��蚝B�m��w[�'䴥˦�}�7����2�3������fˠ����F��s��k�
a�x�ζD�%hH�fJB~�=V����Kɽ�/}��<�@X���W���}\��w�/�U�YR��T��������N�»�&)r����	HHg?���5m/�AqEO�j�{РKa����C��4)��,��L�ڐj)��<z^���r���ǞpM�4��}Cs��)� �{>	X�w�y��\�b�IQ�yb��g�&�<��Tz��,C�,r�O(�b5&i:r�(�uD�3]��=����r��BJK�n4Ue2���ӻ����ti��T���3ܬ��[f+{!/�R3��v�>�l�t�U�aQ)gArs>ښ�j�m-TP�"��v��>::z	��� �q�;��?�_E�au>��(*�!T����\� ˝ޤ8X������<�f�f���F"`lCrJf��E��6g�|���T�F�X�D(9��H�WE�����r�K(j;*a��%�t�3�~�f�I����Q�08Z�0�]�	�	f�kѽ��Ax�]-ϴ;���*��Y}�+Pz�.Zm5�=x���$�Y����K�����x��D7�\��6bad��=��$��R�qg2��0�0 ��6����B��,��v�صO�D�R��#P�WB�5�2B5NIa8�(�h�)�w�c4�:�hW�����fj���舭'r�	�]�! ,$m�	4�(w#T�i�^
�<�H��.�;N�LGP��=`�V!��s@�Aӈ�,{zΎ�����53�,�fp��!��`:���I�W��S�~щ22Ժ��b�PϢ�RvFh�O<��߉@hÛq�Sa�j�L1� =�������=��;�(�t�@9��\>�mB�ौf�.�N��p^�J]��+�B'|�̛7�%d����QY"�<���W�������k�O�.�g���{E����͊%�Z�E�B��8mP�_�<:U�Ǌ	ve�p:zZ����#���
���A��=�����X`72H� k+�B���y�%�����ۊ�$j�U�2���	�v��yڅէPm`���۪g���7�g�vp��3�Zo�V�o��B^|��w�.?�y�l�Þ��z ��ͻc�۞���E���N�Z��b4?Zh�g�L���fBy@8Ci@�+�s��J�L�/�D��u|e㿾��n���WGI������+�N-w@Z���ͫ�d����Ǭ�E��s��!Q����=ǚ���"��
��¨��r&���:�d�*,+�V$�텥���Q��r�M���Et���;��@c�}{(L��2����
��dȷA�W�G�yg�k'5�u��"�V�=5Y�2�"�UZ��b܄��C��=��5D�EY�uMTX�zzW���s��BC�6�@Pz8�,�6��ة�v�����[O�j��4C���̴��g�}*��Y�WQ������+^���K�ar��B��{���2s��m�	�y$����Ybu��U��A�r��c�I��ͼ;Nx�\	J����k�Nd����f|UtTL��l'2�����i�_͢X��0�P�����;��S��A��}�<��aј ��MR����ٺ���;�+������ Q[���8��c��KR_�H�\�� �I�}U��َ8K�) �T��F	�p�gj�d̴�l��糼۰Y5#���� \���gj���FxG�4�QʘTǓ	T<�'��IV	��)u��<ʖn�P&5��͸��SPl	l�"���,KR��3��­�ѵ�l�Ԫ��ƺ��_���ws�w� !7�S~�T�
.���,��>q�i�w�o��QmP����BK�R7����P��@Զׅ�V���)5�@=s�|�Jp��U�M���kJ<Z�ǿn�ʹ��_����R�`�/�/��0��}�%�e4,ۭ>f��&���7"����e�z���0�[�+����\�|P�cA��|dL�$��� ��	��
UI�uG��˱�<qw#e D�'#�fW�<��:8�,,��E�\c�?t���h+����:���ZFu��፻�n��������'B��V8�4tf)� p�v�p�)���I�O Hk��z�|�d<�1hB��Y���-q��VBԜ'����ú�����ZNi�W��r6�+bV�ȵ����+6��@���/���He��!���e%[������#6W��S�Lڒ,��.M$ԟ�0�}c ���*��<�Ր���Q|a��w3^S*��b���8�7�����ӟMJH
l��c�m�"��%!��w隷SU�[<�����^� By*��-�*���唨�EVҖB�Uϗ�h�?��N���<��_S�o��YC3�.�eP-��{ޓ�?ĢK$�-g�:��$N/�PY^�;�;#Y*�7zH�! ���~�3NaiZ���:��6�XT�����՝�8
sY�@���꬇g_$�;V��)�L$&����'��QyvK܁Ӓ�S������T��y�|��k�R
<H�h��96Ɇ��4��Z���yi�Qs�jeZ˔u���4}q�Tn�l��c��2{?�z�)�t��*|���[^���
��N��j��>^��{Ou��Ɂ��j鰈Q�<\:>LT�g!IcR?�'g�M�X�Fq�V~��n�͕��?v�WΆIe�}�!MEd��Q3��"�؆'M���3����5#m�ā�'4ƹ�k"�{ͥJ"T(t�i��Q�?�#$�$�sp3�g����B�6K|��8,���'��;|CY����.�c :�Q���г�?�؋�p�T���!�Ș�=x2-އ:�/��!*����p>�� �����q����G{�-�̻K��Lֈ)m�<��ɓܔV�,��[�f-AV*N,ƞr�� ��W��!��ܟչ6o�HZ�h��$ivE�Ί����ޣ7n�tL������,rH�Ï&@�;2�s��!�޳-���c��k;�3'��9��2h o��Z��[>甯��W)g�Ȭ��8��� �k��[(-��;-]�;�1�7֠HN09��z���IQ�pf" �8%����e��S�Ã��z��B�>�p[C���E��I�J�\9�`���c��M�(1BU��/��I�Hh�� ڙv!:�8����UI2����cJ�Q���NJz᳑�4�F�����A������Ap�1�#P���2c<3m���s͟Я�X��3!��I�*Ъu�BK�VO��F�)\ ��%S���8�G�j�iP���2:QeL��u�.vS��sD�lH��!.���7�o�/�×�Ʌ��7��˸py��P��/�Fh�.��K�X��s�$�8-1�%-�����>�bQ����(��%��gVh�K��9���p�0�,ܴI��O�n�`�9KrGZF\ա�ڦ�疕���V�9���ŷO�R_c��������%Ie�����= XM×1<!�e\Od��>�b�T�)���*8_a9�BYv,Ԯ4�qJ#H��\�ځ5?�j՝`�	wE�C�������ڹ.��+����xs>���IUN�~F�p�X��ĴJ��[lp���,��j�9�w�mdOk�'����ݸ�t��F�K�դ�Ůh1k����E�7ā��]�sJe_"�SZ�N�w��v����q_y͔���7�k���'�%Ŷb��s���b
;�L�e�|�3C�c� #�6�I� 󓰇�]�7&�@�ǚ�c�۬���UaH�{N.�g���eflUDO�!��UH#�;B�?�H� �7��k5C|�Y����
)X�&0����y�|P��=:=�?���\�O�X9�=�"մ��O�[�	�[T6���2J{� l�5��#֢n�qz���.ij�e����i�x9hWƈ����2E�"��RiX��{����{���u�S`�J��J�.��Iyͺ��TB(�ְ�g�J~�:,X83ۻ�6�H5{Ί
�ϔsz��A�S]`�z�뇑r^9���.$�!�<!�����!�х�sM0���͇v,�	�luM��gS�<e�~����\iұ$�����e�s���wr�w����/e��1t���cď£��e��.�1�$�b��T��!��\�/���I�]�74�9��t�&�b�����A	��,⻞m����/��z��������|n�L�����6��	Cw5;���\%��6B&SI&W���u���\�`�k0�mO�\>�Q�:��u��/I�G~��4@��6S��̹n��D�>����\�Y��DD�h�l��4eW:1e��6I�#?� �����|,C /_#=E$�KL�nT���MqeYK*��RN����]�L�?�Ʋ��)����3��:"O��4.Oq�J��!��}���1�A4���J|��)�8�7jq7=���2.�P]l!�0�g�]��U���`L~ߍ��3�����7�F�a�F�>`��s�����]N�w��<K!	��{�ܾ],CA�ዝ��� 0Z��<B9���P�!����_��7�J��KBI�&��7�ԓeث�g��