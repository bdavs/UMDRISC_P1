XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������fPt~�_)c�G�����ہ|D����嬃�/�̰Y�%�Wm���(K���N�m�(+�ڙmn�A�k��e�K!!���4E�Dqx�6��N�ߗ�:��d#�ݠv�Y�r���f:.����b:�%k�N*�`�Cl�U�d�y��5<����B�����e�q<�J�j���q@@l�B�y]���0�>RnW�H��Y1��(�?���k+�|��*�/=/uN��r@8�c`m7@b�,15h��9n��ğI��uK�e���xJ#�����0��
�O(�.����Q~M��*�V'��߸xD���=���q%�KW�3L6z6��x�~`*�M���L��QЋ�e�(*
�)��O*�GHZm�^�0%E���C��u ��S-�k��A�-��\���H�l�@Ҹ�	�,d�H�<'�~`ǏE���qV����������Z�2����u�����kp#!cQ�[@����=��j�9�XX�?btVH"�`�eɍט�N��Տ��:<�#��Da[糦D����cL����IK�=�;����q�Ɋ�V��U
"~��d���j�i�nEO�k��߿�%���e�Ј��g7O�4�D������O�e��6Yz�C����~�`e,����
���t�<��WH&�F"���ؔ���k�� $��I��V�u9[�
��&��H�����<��phi.�Ƶ�ԑ�����S{�� �/��[��U��)bXlxVHYEB    c763    2600#tX����}���SXM�����	�?m��E_壬2Cj �z�F�8l������Ru�Pb6TFS�jm�n�K������-�Ԫ�o��U8����I	d1�jZ������h�Lȧ� l����B��d������q��A�D8���۲��4ϵ��.y!.���ݘ��!��4J�H��zѸ��������Rt�J���4ߏ�bg�{�b�  ���s
	/�<��X/@�t��O35l}�2�nfi�%��R?�]���cО��U��q��q���M�	e|�\�}��ճ"em�J/�F�_� ��k�d�+�؇*�I�
�a?����`7S����j��+xܫy�Qy8��9���}��}��
�\���uNxhz"�[rd�֏U�"`;�M}��RY��ʞ����gGꀭy���ʋ�2�����,Y������Q�繠�t`u{�`+Z�I�ٔ���eR@OA�2�'Q��k8���R�6W���P�2���2��o_y0]�)�io��?(�D�����L|.#u�;[��d�dCp�Ď��O<5@�*�h�1�y5Q�3!���>��_V=,7�{���IP"<
[ZT�&ІK�!�m?�z��$k�7�I��oe�x7,8JY%lw�X϶�t�
7�k5ьc϶���0�r���#��=Jx�X��y���$�R,լ��
�/���6�;����?�9����������h_���no�Ű��'���4��%Y��S��{0���Z'?>��|�F���XX��T��%b��r�c@�~DLj���׺��e�bC��7����ڠ�N�X�����v\�������I�7���ˣ@!hK���m�=��o�މ�i׳8n�+�KǊ�]1���&>L&j�م	��������T�?޽A��ǳKmE�ș$�į�e*��}��q�:It��� ��r1?�Ҹv1�.X�L��3�@��%�9�uo�/����/d��i�{TD��n�����r�2E.{��r��(��}O�\W[��=(o����������Wn�mm�n�.��^�X1��xU�bX�^"2�X?��'H��@a���[$��h�0F1o ;�߉�O޶��Zf.�䟂<�X)�;�GԯVz!�0J�����+	�Fؚ�A�1�`d���\`��Q�P�N��ٟ�KeӄZY.�=D*����I��eHE�.B>s�#��)�H(����l
j�qJ\�#[׀�e�������%���^��ĦeFV	����ѯ�䢢�# �-G��x�Ϗ�v� `t��?�2�ꯑ,�f��EmC����� !�]Oc��c�?t\�#�[	N����iSr���s���*��z����W]�
��\�Fv��v�L�WI#��fk2���+���!�#����mD݂J�c�����QZ*7��g_����M����[�Ms�>�V��G [���W��j��e�&{>e_P��Ǚ�ue�\�Q.4}۷i��N@3�g�O����̼�@��Ғo�(=뜯��sK��u_����q�Hp� m��!�g�6����9��/̀�|ˊ)W@M�z��d�3A��Z+�_�}�a�-���?!>��k�f;���u#�(tz��N3:��2��];��H۱��Q������y*�@�;�9 �iF<��Lv&���h�C��4Y��.�̟�׫�3���A��c�h�` W>Ɗ���Qe�����me��?��f:�)@_v{�Iڴ��tx��uYA �$�n�uE��<�3AWc�@�"����z'+`�Ae��C^p
�r�� eD�������ZTe�X��e���hR�~8��+f�+��Jq-�� Й��7b�H@���<w�$</��L���du)��Zz+�svƏ�Y-v��mts����l5|5���tZ���]�l�jDW�5�a*��Ð�*2>����y3?��L� ��oj!�����6xN�C���,��4}���4�;��	�~��91�݇��w���Sk�F%�[��Z��Ad�JL�cvJR����9�'���e��\y������x{���,�E"��X$H씴@
�u;/K {�+�Ͻ6�}�cf����V�&�ERq������vڂj�9��������F?�7J��0c~G�� �[��2��9X�2"F=�f<|��nl����9B�n��-�jg]�'�#�ќ��⮷��v�L���h�}*��Q��q�r�+	��S�p��(6a��gyEo4r̟>c�v�ଅ����'��\JZ�Y\���.�v��Z�@e��K�4˧�;=q�HU�k�g`]3��J���$��O��}�A��p�������R.X��̬�qw�mAj.
B7��������a�*�)NP;=y�$�q�	�"�j"��f,�l�w*���Ky;\^c�Y���ym�����i�Y]�g�`(j�Mc}�q��l����aMT�/zK��fy���Q�z�U�ݸVg�y�	N�
��SX��-��JR���m@�����n-����&�"��[[|>5Kp�U/�2<d��w�q�O��u�WE���a���hھ@�I�Z��⋆U�3u��]�� �BeWU(�a:��Rkr̓���Ʊ�����Q)KOLIPe���->���&FL���<,w�Z�L��i�Z���¿�Źa3����iK	a�߮��{)	�f�]�UG���˜��]n��3ף>X(���/��N�d5�Z��	{����D(
w�v�a=�X��j���R<���ds��P��kYߪ����xQ�]����űk%�ƴ���9�8r{|v|6�J�]��3a�"cTkLidݏ�1_J��:4�!B4�Ia)���om��`_&��~PL�h&��k�"n�U=r�F�/67N[j�ݡp��qM-8
������������ �q���D�ٲG޻�o��*�ƛsG��a�s_�#*�"�����)���Kul|���4�]��;�CE!�E����f��L��O�oEs�!땫Y�\~�g�>�A��dP��+����<�  �]~9+#�X���-P�q��2i��@>�s�`,=OgD>�ϩǸ��3�֔8u������2����[DOM�,����o���){.-��W� l�f��㘰zyH�ۄ�����GdR0	Xk�#��89nsa��AS�� h=-��d#it��Q�wXVuxc�[h��П|[������B�x��������$�x�y�1'��+����	�����,�t)���rp���Y�̅тC��"�E��'�z|r������͉a-D�a�
��~"�UR�8B�^�X{"�_1�KUc�p��߯S��|jE�Z�H�IgC�!:@�R�܃�'���hj�
�i�&O���̀ޗ<w����)@ٓ�x��|�B;�t%�F��4��kEo�Y�� o����󏚆�������ce�ގ���}�n������^�7\�%�������K�d���tz�.`6Ql������,<j�WP����K�O�8m�M���cQ�7d� l���@'R�e+J%�� �R>�k�Hh�T�F<����T�@؜'�#��:�฼U��=}�0	�<%a5��u..	���n9'/v�v� �s��Tᶐ#*����%�z���/��Bc�b�C�.Ak��=��˃�kpGiz����;'��y�AsgZo���mf����j�_+�i1S#��,����b�>Hc�
7N[_TϛT�u~�`��}a a�S��Hw�=�Ai�hO	C�`mF� xwj60�k��M��Q�������F�>��v����R$��l�]��̜%FU��4=��ʀ�ޒ�}ʥ�[%�`�\��xS�(�c哙��ќ��)�D��Xp�ub�R�F�dp��*�x�P��y+�t.O�F~W������M;�+"? >�q�~b��x��8f�\}�t%�Π#q����r���Ŷ�<0D�+%��������T�i���߫����s=d�+7�,�/fb� (zz�Ʀǳ��t��1��6n����L@y*C�X�UP
y��D�,ψ��9�#�.�H�� 8o�ִ1��a	p�D� a�-�d����1�'��](����@wGo�?���	���/qV���qYK�BN���P���uA�-t7~h]��������2D4�vT?(��͙k)�8�W��:�KK��#)�+e�*�\i���&ӭ���V�A$�5!�僃Q��+kb�ף�A_Ug��յ�'���� k�w
&Y�l@i_�e���uI���Q�Q"���`���pKK���yH�qm��3��G�A 4(y�LL�l��"���Ӻ/�ך�� �^�<��bX�
~���m�1Dŵ����52f[�nǐ���
yw�1���a��]v��M2���K��Ω�	���qzr���� ��o6\�2F����0��Df����g׳�԰��[@�6^���}�"��5��{(W�3�ԃ7�7��{��|^uX����ʗ`=������⣔�W!%_g[ƥ8\���y�FP�OB��Q�7�ˌ�����Au%d*3�e|{�oL�(��=�᯴4nXs�HK�Ru��*vqL�Lӆ��[�=/��e+aw0��_aģu�LBY�Wq>����:�4ũ+8au�����6��t`�@E\f�����C�	�E�ȏH���C���_a�����ٌ��H���ng�&1�@a��~.�Pq)X��'UU+�S�ݬ�KHНϷ���"�B�f�q��+֚�SQ��x��((� �Y�g[�w#g�}w~����^���+y�k�Q e��z�����`,���骹���	d¤�H)V�o�O�rg��Z�����o������gLuk���|��q#�U�=��Az�pAsy?V�r��&���W.�t��z��?ע�L=Z<�Ao�-��p��껗���^�����%�$fG��]��N��=b��ީb��Ń��[�P*`]�S�6\8V��E�+���$��NM�/pb)��"b��3�V��`~���R�0�G��z�>�׽|��o�޵]���x���_����e�fr�=��jޤ:~%��]�7�/�&i�h9�J�O��>�@�����5�J5j������[n� ��Ʌ����w�Z �0}M.%��
|(��(�ި�f***��m_�Ϝ��_���٭�ba��;+{�n�a�N7��2.�v� R�P�1yc4�2X������jI�,̂�4��{����»��QbU9��e��J��[6o5q�J�?�>�3�3�cp������X�j_�~����r�q�����4狍�7x�x] �o`�?��C@����F����q{~[&� �P���֎ |�k���[�Q����S�eAz��
�n�����/Ծ���b䛑\R���.������Ɔ�[-��>�ǆ���r:�>.V�(�΁o|��e.�~SsYܠ�4���<"!!_��$�N5�>����/��.��J���R�-,9L�^��9c��̒T���S�"�ݤ�?]q�<�&�|/@�[�*7X��|�a�3�-�%�_�:��J�qvWL��(+9{P�$�VՎ#
��7_��lzKcw���ɗ�5HiB�!�xz�6� �]�$�gun��y96�?�^�N��ِ�g����N槈��H�!�	��2	u����(,mRM]��%n�g�1�?T�qFn&���� �����L'~�-���ɕ��&�Ŷ�3���.<𽯻��_bOq��%j�A�lckA��1�CB���:����J�N��(EWv��<��
[>'�c�P#c��5�0�P��0��w��sL`*�~U/T�y���G�"Q����qJ�ꉺ�9��U���IIP�TqI�gmG���j�.A^�I�$�Rւ�[��%���	y��V���5����������U�l���1�ի��u/�9�^w�^� n�(t$S��eF"��0l	f���I�o1[����w�s80$��}���k�#LXM�|�(w<�cX�cf��;ۭ��T4�+�q�z��űsA(Hv�{7l�e�GoJI(�Og���ϝ՘6� ����p��v�e0���z�����U����>f"s$�yȡ��9i)2_2cV7Q�������V�:�:^4�\E�},�>?�,�3��%�5��=oZ���+��no�C�~��N�g��)��!���y]��Og�S|M�'�/qw@�u�����D@���궖���6��S1
4�v�`�=��S�ͱ2�Mּ�����h"�LKG`=	�Ղ>񆮀�E酒)VD�� �Deʸ�V*ϛ^���pjY���?�!|���.d��6��j��J.�n��wD�"dg��n����{L�a�����O����ID]���G-cp�W3
�-��l_�{v���@��B�F�[��GoU�3Ҟ��:E@��-�%K����2����!���N,�}�����^U z��9q��o./^U�v�S�g���9b�@��(ҵ�s�4���bU^�!�����c�J!�Uxܥ�=�ȳ퇠�#���Y�]���Q1c��w�N!>ht�ݣ�iW��q~	U��wx�Rh����uj��b�W<7�+F��4&�|���6c��g7��	��)3�Q1��vun�oERE|T~�YT��FH�cK#ƞL:�����G��R}S�/��T��ޚ�.�N��f�%Hة���Y ظ�ݦ�C�U��}�T���N�(-��	����\&���z��r��<H:��4/���P�d�@�Hn��czw�U�%��~�������m8«�#��lVT�4Ez�t���} ��J�~%2��b_�D��\��$�,�GS)���N����q��UO)� d�C�*.����U��Z����I�,��Y1H
a�e���cΙS@���8���CK%�ץ%�e� @�0���\+�%��������[#�`	h^E��Vc����)���5�@�UfJ�Hv��k���A�I�ź�4���aG����˗4�7(�[��Q,�HTy��>xb�Z$,W���!��B�v��P����_-n��  ��w��p�(�?���#r�כk�;�6fUM�^�d#*��ւ����Fv��6A��>�2mi2�L�������y� �'rZ�Η��TT9(:�)l=
���Q;���y�i{D��"Et��N��IԳ���/���ΐ���~�A���(j�1$��au���s e8D��M������1I����H�7J���0��r� ������A�&��x+=e���^G�h��Em�g���~צe��5m�c H*_�3�����螛��'�_0�>k]/M,b��N�]˸aǪ�V�
LN���~�YԭF�ѩ�^3t"Y��P����T@=�~Ŵ':����f&�lQ�,���"���x�s8���C�R/D��0���Ҁ��;�0n��B���'���7�:_����!m�52���1s�)\�����A�.�`c$���ŧ�l��X'�D�HR�"���^��:وJ���'�J�s֬�:��ץd�;��Q���\�@ց�kj�,�z|��ThѮV"�4��"DR���0�挴����2=mB �Q��z�V�b�0��R���D\��y�'��k�6��uD�'��W�h.��Kf[ِ�Pg!0!r���b5����>#1��n}hUz��%����Jv?���7ܐZ `�3�b3:�<����"G�����S �f����S}�Ax}�V����?a���b.!��d�Ӓ�u{y�����ׄ���{�J��4��_�P��>��Y2IAO��������)B�ʁ9\����oB~�Y���%�=�U���>������?c���t�ujv\�o�������kJ D"D�'EV�{��fXHO�����B�+�
��W%l��5	�z��0S�T��I����>�w���fY�ě� kJ=���>��Y���)C}r�I���57���K龶���k�}�%I������i��F���������ۼX�n@M���?��x�.��\Iph<=����OJ��g7��K�L�[s2^��ٚr���E�\��bi��J!z73Y�h8�,D'��s+1��c;	�I��U�׼5qK�`�[���S��1��A�WG	䍅��|�l֊#�]s��-�k��˻��n"��֔�R��K��?H���k��F�!�D.����$y�vZ���S*UM}�ƴ�m�L�3�ux@�Q���3`�W�R�t�ϐ�;�b5�x�IN�{�,�_��j�PЬWg�-H_޺�S��7%�]Q�@#,�s�<��ʷ�5ўg�3�,��2}c`5Oe�w�����s�K�#u����ە�0�̊��V.Y:/Y��]�܁C���j\踍x�G8l�Xc2��]�Z<-��؀�1U�ҠÒ^��@v�+KuSf�������$Syw�0/|�x�sW	Z��X�P�c,����<I긦b�*:8���
9n�:� |j��ɴH纎�3�J*���d"��T��5c��Acw?����Z#�$��A�A�bEK�&��E�������Vh‹'�2N�_{$�P����C�EL�}*�{�1�4F����Q��4�~���;��^�����)��i�*dN|ڍ��f��p���ض���,���Ƃ= ��W�����Z�˓�b"\Jݢ$H��L��]:i�7N�d>T�}�Eq��V=*sp�1�h�F�&�mEh���7��ɰ���tF2��L�Vɶ��JL�����=r�mX��F+����om[�}V�x��^�ڔ�Q���(�b���e5J����O��g��x̑��ь�po��oF���?b呩��B���I���[�8�\�T�J��mN��#�����Llκ�X�G*>h�|��:Չ�Dm���v�b����i�!Y]���^R�;�>�|"&�i_{��^x����K�����7.� 7_9u=��UC9�FjU_���:	�$� I��gܰ��HfG���2��~�_�l��X�.�P���9��ޢO6��AT���PK��M��h�+n����$���ÿ�5��h�(�K���p��!�.mV��:�E�qA��N�|���]����g�c.��l<�,v�d.Wt�'��������$ ֑�"?L����}(Lr����T���ˈ3��!��q Us�g��;y�)&Q��'3�,���(j]������(����T����F+�"����%!��$tǲ����1hm�Ɵ(��Ś-�Xsv���V����A����,���@��dB����6��1�$b��}-���t0ѻ�*qA�����ƿu�Τ!yګ:���������]R�����:��|�d<W��!��b8|o�)$���2���wQ��&(·��%��� ���WW㔦K�.�N8�l�����i�Al:z-���w/�5��a�Y��rF�=u�[D�-1�R�%-Ҟ�@"��X�H�