XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�ب�,C޳���e��#�S'�o��faZ,:��7��gN��^�Ç��[���F�UE���)��g����݉�?r?$Ov�M#)�vɝ�P�MsW{���7=_����/�8�*�
�:\�]u�5�g��̇ �wMF&��:�\��鴊[��D =�R�)j�^fZ���]���{����Q�9}�o��\��I%�gz�̪e�];�r�2���]N�.����8o�>�N )�|8�s����N^�ce�%}Z�P���O�ii�B��%�<HU8D͎x�l8��J�[㊢t/��(c3
c6E&���g+���C£h=X�B��];�1k
74�S:eg뙦��V�@��p����D+kbq�N�����,pښ�v�AGo��%�,�ܙq�f�㭼�B����np!�hd�VP�P���cD�;s��Hk�:qI�#��BY���@�ɻ�H"c�����G��G�r>���Nz&6��È���t͌�㤯 ����қMa|�+�1�Y��լ��^�$�"_�����c���&�R&\(��ߢ@�Vк}M�n�w��O/�R��8��;��<=�A�`�+A�0{/��%�ny�^yI]j+;\����9��X0+���*Wo�'�5�"ԜZ�Bv��ƜĬ��z�x�Eeoxs����Px�B�T�:d�1*i�[5���s����������BFf��T��}����#�d���5]`����Jb�M˭�@%$���0�vrXlxVHYEB    fa00    2560�S����1oEx��~yis�WT�3��}�sNO:9�P����u���ɘ�{��P�d�-)6��FǙX��7��X>����+�tVk�M��鿆[hc�xqz#s�!��T�%�盼T���)NG"�7���)���N��	�7��ym/~���Q830^�oόLΞW�_��Vn�K���I���lq$u�V�.��=XT��_&<��Cn��� Cr\'�����}00vb��O�����FG�d�'�7���Rs��ˠ��m��Ď:���G�W�.x`�㉅&Z��OI��t�kN"n���U����m��9(��{�������P9\?��N43;�����+F�`}�k��_o�9�O��«�+\AU����׋_�iY��O��Ż��J}��L(�o����MźM~_؁/<�ſ�gܝn��Yߗ"�z9;���훫�0.	}YL�	#Q7Yڃ
_6�8��¼�ٍ: �i�z렆Mv{�qR��҈��TGuY!�z�S	`[$����ks2�|#���O��lx[�#��?�1}������3�OD��:UZ�Ì]�u����籷(���K�v�uO�*��T����s��"rKR酛?�7Kd�4��: �o�b�����xpT�97J���K%��^s.0�c(��o��x��k���'̔����w�	4j�YhYR�\1sB\ZC#c��_�t|9��a�E����A�&�ғ�=���}���[������w�[%[��S�O�@I�G��1����m��KAeWX��IlK�2�j�䔱&�,�E�_Jo:�H���
c���P 7;�;} �*��v�9��ۈ7����5u���u���,u_9�;I6W�5�7#�+,|^���z:D1�	ϗ��}�m��ߔn�[�����,g������4�~��6� ��8G3�#���z�2}�Z隹�O�T�&��6��M%sK��(���-b�g����2�t-�����7���"խ�l�0�ƪ��Q��DW���)��0��#[ۍ�'F�[,�h(25D@K��i��@6�;&��h��������3y�OF�A>���I��ʏ�����a��HI�
<��
�\�*�h��4~�J�@��ƉCAa���/��ƕ�U$��K�����H
��+�Y�#�HJI�"�%�#æ.$c*ҟ�8�O9�)4E�شk�r����A�n��"���H�ce�ǂ#�G)*ݧ��<r�T�����>����7t|�$w�v���n�v� 57j�ߦ��ZS�˒�YȢ��G��5���<-g�*l����~9�0[�>���v2��4Du��eןESRKK�y�T3�'�ha�N~1̆�xL�o=�XJ�f��Yx�1ڧm�����lлf�u�f������B�@�?Rʢ�RA�P�L׏��������N�ӄ2�4˞$A�w�_iu����k:#L��i�t��d���������#{f$P�yp�Fz�뜯ˈ�c ?�\��
�z�P*��������;�7�t�����(��SޞU�K|������QV����"ĝ��]�R�#�Do����jE�;\hqt^���%S�`w�,�U���O�1��]B��yJ.�Xx+�ϲ��.�y�P%���- EDF#�1���F��3�T[���7��
���)���p����?�{ $��g�pg���d2zN�赎՘�J�{{1��B�S�ϒ"��_{+QoR������u��1+9�Cs�b��kҨt-��
��4;u#��l�@o��]W;q=�IZ4���}���P~�o;��ԫULiM���M �ʋ���R�r&n����(�M���K6Ц:P��%h�<:>�� �[Ц�6m��吔�~�e]:��g/��B�cH��͡L��@�f��C��:�sC#���!J�B����������tFϦ�>Fx�P��4��ؓg<.Kg��ɶ�(�#˸>�|����\�������?���f�&��o�:�6)������(4���;��9��`]^�/������J�B�+�p�a}��RD���3?6K�)�\���q�gpH�kKM�?LRpR�~��0n�"K�E[��B6�-�*��@$�戯%��<�0�������)��U���@��wf��Ջ�T2����l�5��H�r�H<I)�z���EX���������,�KO�A���7��'Cj����	�T7���##Z�~��/ͯ�6��l�{�ۑ�i� �TGZ@[����9��K:/�
�)�����H*��s!mE-�ԍ�5�q)h�4 �U��^ѕ�+�$G�u�x��>���?�j��5@Y0���ޖ��FOw���\�V�ٱjGtU�CL�;5(��6�6֣�$� j=qBd͹�������q�);��W����C�u� <=�"�\&����Sݡt� GPro'2��h��0�9�Z��;$x����a5Y�Y�"	oŐG]KL�tX޽�r������-P���ƨ����<i��#p��6��5���Ͻ�=����O�Z��o�@K����*?L�[*���4����4�
2�k�B���5Bː��1��\^n�57����7˭�l^u�k�G����3Jk�����ږ�0� 1-��a)�K}w�@`��"�<�>��9?Ǟ�6�RDCl)_�s�8�p�Ɩ' ��&a�Ȫ�k�แ �Q1�[y˧�˴�6/o����*�qu�e�|wї\5��G
o��~���GSW�N�ë��AOQ���C��O<"�yl,]-P'(����5C��b���]3pz��_#S^��|���C�`�Y��̰����5��ټ���ߋؖ��M�CC�։l����hO���=�-�s+�R��#�|���q~�MͽH>γ�����G����M��G���G���60�H09�Ȓ}K��L����'Fu�)��S���l�U�'	:_�D:^�"K��u�*JSˑ�Y��X/��N;F�����T�ǉ!�bbd�5�J��P�Xp⒵��� ђ�6,3��f�m(���!Lex��pD��a��w���n筒B�hg��W˞�U��V?�$p�o����@���g��x���8i�����9�!���U�+'�uDa�� Q�;Es3�K���J�6Ϋ��ˢ�U8]t1ژZ�?䨽��w�m���,mP�z5+�𕪧Z���������\xz��=��߱�Chl������/W��jCqyh���h�z��ق~��෻�>��X�E���f��G�:�و~Txp	>�|'Nj��#���4$�Y�q��B-�o o�Z���Mƨ\����X}hov�"OrW@	u�l�#e7_�"��ոɡ��m؊��D�c:�#�<�7���ϙ�S;��Y�}n�ǌ�]��S�9�S��o�m�${�>�;��t��1Oi��2�D���Ġ��������b��%����o\~���tK��_��>��1v�\�+�����E�9��]���L���'��n�覵��:��a7��脁�����O ���Ն�i4�~��d$���F�L\p8U��잾�2�F2��H)���f|�����[��ћ�{�ʰ�Sr�ZA=M�ta�]Pt��[Z��zc��H���1��V[�N�f(�c	�/�W�t���k���m��5Aj6����#ݳ�����$N�1��7[��Z���r��j�0���I/2�Z���xE�V�4�\@�!,L�A���=��^���(Xz�r�~}Y�r���0�.���zP��/a}�*�z�i�>����Cv�1�q�����Ɗ�T[ �g�z�]RjQ/�����e�R�ݏ �
��0�h/��)ڭ�L�[梼9Q�+�f��� �4�m�5�@(jg+05�A0��-8����>V�PܿLf34�(5 (���T:������2d5�L�F�}�۾[wͮ�lF�٭�6Y�CI�1� ���ӓ��sa�$Υ[ۤ��С���������J?c�F�B�rQ�#��i:� ".��-���l��)#U�7e�0�Imֱ�H����|0�_�s�/�9�粬|�k�OE`F�_t_�Ơ�Y1˝�È$T�y@� ޠ�]�J�+�e�JX�ҵ��f�ue}�X��[{�sk��dm�x^u�j�;P£0ɜ��Ʀ�:XH!�O�
mfk�!�a�o"��y �(�=���h>j�C����ME��(D\�� ����2]`e�*��ҒKN\�綄�:q׽t(pX��e88q�k�5��|��,`>�	��>-�Y��4��K}Mt�a'���#l�5��l'\�n���DI���*���y�8IU\���7�5����h��E{r�,���/�2��l7w���B5<�C�"�+V"5���&J�Ԝ�a���_O}�������ASw��O�XJ�
����F�A���*-�J�Ƚ��z晝��⹼��ax�rj��N�.krvx��8����ܨ\�)��b�I;�^�	��M��7-Ϋ �#ӛ�d��?3H��h
�3�G�y2s��5B�"����Ű��s�
;�6x�<��f�ȁL��+�F�3��*�6*�����CBS<�����4K��)��[��*�"��[�n����#D��[��c�r���ZM�?�^�A��St{An�Ph�0��-%���@ɿ�\nyZ������s�yy�W�Łgpy����Q�iDp��v�KdI�<�NZ(��$����"}G~�$�������1��+~Z��V`�oe�s��U�����_hC��dB��tD��|�ڥ�+���=
AĪ:w�N:�vL�]��c�7-��У���rM���k�lŕ�ߎ֙ο�nf�r��s5��VΕK� Xc�=��?Ul:`��$>��ۧۜ�ӑu
O���]�-��������?8J�1��_�4W�OU�{T#��(�Pئ®��o�(������P�'��W�*o� �����r��gC�'q�(���Ij*���sC��g�����Iqb
a�*�˛+i&k�^�X���Sb�� �E3��o�:�/e/8���$\G��������U�=��p")-"3�0(N�S;.S�_�O��l�fN�1��:E���Q"��"�d�c�5��ъe``���IP&�IX:?�m�>�f;Y3���t���A5��ȫNY*j�*uZ��p�b�oj����,
���r��~�Ei��:�00?h#����]�,W�O4 �Q �	��j_w���ϋ#��0��`�B��D9fЋ|�����H��I��~�����WS�
/�td�g�/ƞâ���W�W�I_`���C�y��w5_�PX�^��P��h�UC�|�S�2��	��j��7&������mh����։���]����W@x2+�r(�k;o�<�80��Yӂ*���ՙC6�;���Љ h2q�z��dr�)� F�S������e2[-M���hKΰ�zA�%���IT�y���!=G�?���w�6qUW�m���-^��@��|9�����L�Z�0�"��#ⴏ�ab.gO����x��չ".�%gWC;&#��&���\u<�AUA��䅈�L��OԾ=�T�Y�|��2�n���O���@�a��*fYA��d�W��/����W�eC\�O�i{��|�e��/�h��6߈�̀	�k����@{-��H��t-)e����u����j��VD���0G�V!G�̼�� 8c������]��[��+jN~x��4���!�w�5{{�f3�Fy�b>zbֶmW�Q}��ʼd����F��i&E>2g�v ��2�3�U���2j>�"?�Z���VE�������%�d�*n$�ud-��TW��B���a��6�Ҽ�A��X�  ՝(�d�CY���z\
��1�B�<_ >E�z�_�sUD]���A�ù�X�`�0�K~ZB���'��zw>&2N���6�$㰚&�_kv�c��u�������S�*��	7��P��o�<"��D��Hɥ7�Jz���~=GW�β=#�̈́��Xln�1f)EsW�� �lk�����m t#�/��
�J؏6�6�%b�	�Ӿ�Q�5�Y�xAQ�f��f%�S�����m�����5-�yt�bO���� :�wJ��XzJ�9���Pe�:V�@���-]Ì a�G%Q/u	?�2I�C�d��;��_�jeHB�U�I�?d����p��"5�s
r���uI�޻Jjc�
�UE��x����8io?H$��|�%X��d��FK_�6��Z���vF�э:�u-m�Ѐ��CF� ����z���X � @���@oS�����e���G��,�Ԁ=������r������	M�L�31j 4����E�M��NF��C���X�� ���!�r�)��*#��.@5�*2�g��z�\���b�^�!��H��B*o��e�� �>^S
�q����Q�p�LBhk�?��5�P`z���U�am�L��ÍPJ��
\��-9G�#_ٶ<6#�8+ÿ�h��R���B��6o�)��*pDD70�_���˯9��0�G�K�j6}�%p�e^�_6���Jgj��G�.�1oh��[U�j�i����DHإ��w�����|��c�Q���=';�(A���C��򕋽3T��|P,�_@@��}s�L!c������%QM�{<��ɜ�*�&��:�zQ���29<�xJ:��s W���h!Gu����A�
�}�˽w��d��^M��)��Pf�n�y�XK�����em�Aϑ��X��%@�v�\^��ؓ+����@���d'<��/׷(L��v �¬u��H&I�|��6���NS�*7��1�x��C ' �i��a�����F&=
�W8�{�>pio���kw�ޤЊ<_bnￃ�݀J9JTz��ɭ��'%��:�w����e�a������'+&4#�<���o��� �u�6� +� �NL�#�����r����{)J���&�ڎEe���hZ8�;�ehu�X'"`��ng#?H2w��c��s����5(ﭵ�a�L�~����"]�K��xk�:�^Pz�رT�.���؅�Tenl�6AG��2��o��텂WP�%D��l���l����
o��ͨ�B��q.:>I+f�K��G���Jl�ѳ�zxI^�H+�T�K�* B�u��0��F'��j��QNl��q� /�����O �̢��q�fW	L����~�lΔ�8������q�f 5e�c���%I��2~���'��o�0ލ�P�h��ړ���'&|��<��f�bЁf�ڭ<����e��O�������Q�#�`��
�R�m�iH;Z�+���n��=�q��<�ڲ�X͹lC���Wd3/�¢�0�Ck ��[�h/�.c=� b�_W^7�	����N#��_w�����`07(r�F�(�ews���EOoi�j�ޱP��Wj��x�Q"c6o[�M$;
�"�U�����tk5�}N3�<_]ѫ>=k"��oB��Byݦ ��Gͽ�^W����Q�mq�H%KT��-�z��J��3{�m�Bd�,)M��6�{�Zp=U��if�	]�y�\�-)F�OF��s}K&���a8�[R�V�E��c�����RW��L�E�p��j�iZ�ZӖ>()&ײ68����{G4�Y{[㔹�-��Y��J{���l�aI��b}O���Q�A�]��:NG?��I���\#xַ������4�U����}�L1AdWB�5��:Z������Rx��X��ƶ�ֻi���b�\�t�"A�$0W�ˣc3��ҎA���g�+���	S�g��;q�I��ᐃ����/%�q5��Iy)�lP�_|��-�^��KU)��/��;,&x�g��]��p�i�$�)]sOر�;���p�o�G����^�W4�y���
���<�i�f�wDL, ��"Z��q9�09w��x�Ce
�n~M��%}Y<s��Bk�<^�Ӕ��IX)xUΘ}2�[Q�B��'���X<&��/c����BM�i){!ϊ���haܷے<�Ri���[�)%å���pĕ�T�(��� m�l���}Î���d�(>�U���<�_,�8cl������%yR����"ߗI�.u���lo�_�/V�y?��Xb����tl���4�
8u�{��������n��2G�|n�����iL��="wޚ��Κ��2="�uX|{C�#:ܚa��K��v��q�C�˔cw6v��?I�~|�䵒k-1��V2�N׮T8��	��Xj�����[�V��V 
��Д��>m1�[o ��Pi���
zQ�B[�Z��詏�ע0J5�"��C�U&�Cx׾����ǻ�t��;�%�z�����7���*���*SZ�E�(�KJ6�adV�S*�t�#Hs��C�C���=��?#fbς�H���ӿ��T�*���
e��ЄVJ���p"�-��E��O͞m�Gr��3��>��؊/�(�hN�?ͭ
.`i�@�H�<�{4>&���r��&�NW�+~7�!u���ZpYn��O��1$��·����c��	��5�ՀK:F��2��	}M%mz��wiD֙�;��K+�Q��9���e1"�<�^����iHo��ᇚ~E.�ƨ1.Bм-����Q�7d��R��>���������FPչ�/q��th��@sq��v9x�W}����2|�l8-�R=g�u-xN��Si>��r�`��g;t?�����/��L�j�x���]���o����8�Y�����8���7�W�Z͊M��Nu���IC�<k�yW5C�[���j7�g(?��H���t���U�uXI�� �Ӂ�.=R��b5!0����c�t��.ם�J�cʗ)Sx��d�v�Wxҧ@�����Λ����b���t`G��|�쪤v!��W:�1���n����u&%o.�����ޖ��:2��߅^<�j�wuwCva����*���(��Ы���*�m(2�DԳ��b����k�m��|�	���}c��"���G�������LÝz1~�~�WyB9G�ݟ�p���]d�����w� ��32����5�2���s��x '=l��Dx'rQvH�ݏ���	섔��R)p�_0ץ!����٨��o([%r��k�Ѥ��Й�j{�,�������D������eEN��+�d���S���8F�������3��B_�/C��{�,k�ϺO�/�l�&9o� �Ӯܧ����c��
�T�p��j��v5%��x��~��@�^Nj���g�3~>|��i��VJ��D�^�A�M|H�����b��_�����2�`��l�����	Ǧ��c&\�ӕ[]K�k�u\�1Fȩ��轩D���
�"	 Jf'f�1�4
hӝ�$��xƭ��Kd*�$�XlxVHYEB    fa00    14b0�^�TD��z��w<�Cm�R��í��H�|YU��G
�����c!���e)�S5P�~v
T�#��-H�+��E���J��������cz�o��S�3�d0@������V�:�iH�y��y �l���edH�a�G�S�'И��Y�ɡ�������b�=1���,h'�V�<h8VnSO�/n\����w�����L��ΰ$-�|>{�D�O��0��F�+�r_�C�/(���(�ff�8K%bǝ[<q�.�����+�C�b�v�^h�/�ZX�J� �m��L�!%�>4�E#��Jߤ��] (ﴫ��/}`��諐��I	*�S���#0.�F@%��#�⧥�:0v�	1�B�#���)���;?ͷ��ڎf\�[I�Ԝ� obr���r00�g:QWI������7��1�-
��oc��71�ڟQ��|؜z��M8��ك�`��^��R;��%t	!����v����I�@��������:-���q��2ei��1����mk�˻��H����3����]�P�`�C��SU���r�A0��x���;�K��38�������H-|��V�2U�:��,[��;_gr��vC�ܼ#��X��`�n*-��JU'p�c^I�4�r�����������A{����Y�Au��6{+B0��\�|g�:�ŗ����NNTpt�n�\-9�;�riJ���ёB�� �|�F������"-��8��ߟ��kP����p�����G�7�/7����h���a�f�kji�P�l(����|�����N�C�������c&^xS�7��SR:"k�Dw�ɢ�����Â'̍ʉ�n�2c��#��t�]�b2��8V=�u�����1']d��_.b���W���9쩚����&�)s4�O3FpنSyN��*�������⿸�N�c)�G�;{k/�B;�< �?���`SS���u|h����k�tL��4�.2�0���=�֕~��RΣ#T֭���Z#GU �,��l%\�&�I��6��듫u���Σ[J�g &t�8�?��(����W\���G ��m)�<�Ny�;�|c[-ĺbW��7Z�%n���Ҋ�h�ʐ�k*�o{�Y�G`�	~�az9���1�1�������54�"Qc|+�4Z�e΀�=��7��z����d����
׼T���e&�o�aZ���^Ϸ�*d�̷���g24>�P/Nd{���Q����\���]�:}SFu���?MdN� �R!������@�w�Y���TC���o��R{)���y��|�v�(��IԳ��B�|�aPd����0�~������R�G'�ͱ�#�u���W^5�Dr�z������:w	~+�Ϝ�����8�qUO����DG��{�EU+��b [������WG�U�8��K�`������]2%�#��`�
̂h)�wp��_� �8�W�%uXƀo�������]Pį���晄0�.(�����P'S�=�u�� q7E|,:B<yG�� �V#A���P��7�m��C�0�����Q�<���}mmǖl�J�-�A�x�~�Ȓ�����B���-U��v�5k�7W��)x�֖�ߤ��I���̻Oeg�`���:DF�nZŏl �>�Љ3�Xj�ǸQ�����V�Ņ�f������+-[���if/���-\�ś}X�&��{�ׄ�� �a RZ���Ό���+�N�<�3���R�٣�GN°�^R�3j�W�y��@h��h�7��#}���>��8�3e��UP�&WɄۮ�u�ɵ�:r8��{ݕ��T�1 b�k������{���I�QJ��xY ����M�l�7#�����HD�+SՋ68���M���+#��Zo]�D+�y��J�t��_��}s-��0ǂ0���q.s�a�%�(�@�h��qZհ �rQ��������o����
f�����������5إ�ǁ�s�����r�?�6Z\ٝ)Ih��$�^�}Pm���w�(ڎ�4:��/-��aH��J�@���[k@�L�k�U�Ar��0^��eZY��v�R���,���qI��%b�8�����L�7Uz�+�>�٦8��~?ə���B��CX?n+�d�3�䠺O�X��-q�а�h>�5�<�X�ٚN(����58t�ӗ�E��a�<ϼV8甽mP��6>� S­vz�v|���{��v�T�7tp9/}�\�G�ϘAh#]��K�5�����l�dt�UI�ʱ�߮+Z��mN�E�>�.6�̟�h�q��vw?a���vj+��҃�b�S&�nr}��;�2�k����cC�Zv���=�prᖉ�|؏�����*����q�D�Ԉǔ<���/��&��1�����k|�9����.VHs�y�bD��6�6!���jW���Z@��_'�H0��k^�@�L�2Y����R^��!l�_�&�M��[{�O���=V��j���=kf�B����+�J��#��IѰw*]�i�����g�x��6O���8-��}BZ���!��d�N10%v���8WC|�蚚W 1BMr�<��^�&�0��>���X�F���a�qt(\���C�,�,!~�1U��?���V�P/o�eJ>oT܏C�/-�V�E�>��,�]�d���,�W�\2@�X��&v�(�j(�%��0��;�2_/�s�����a���7�'7�t�.9����^�tL�\e�!���ė7 �R�r9YN��m��C�6Vg����$��°@�>�
��#ȔX6`0���,��3��W�ߖ�:���s�:�`�R"q�+�Zəa�\� ���{b3�z�ˤ̀�_O�Q3n���:w��|
��?���t����ho7��5��/f+�F��ԓUzfK�H����>��!�&��U+��gr�i���y|�a���_���<�(=韹(��U��fq���uk�h5��х��"eR?1�Ǫ~��^�a�D�C���th$��^V�*��8�_6�*�bQ�щ��I��u���O�$�c�ܾ;6x7{�z�!9��A�.!�����oָ�=���^6v-%���)Q��̹tl.�1ϑ��;�)����L3hv~;s��Q�=1f\�M�r���D��p�Z�NK��P�=L�]Y��Y5Q�y��Fy�o�$-����r@\%t$�-w$z �X���]-���PTq�Ƨ#�L�˂�^���X�w9D��Ҕ��V��qS�$ _9�@c�� �@�c u!,��e�BJ9����j~���h����,����X� �k��R�O?>:�wctv7�Y�*�d|e ����,	��2#��G�7.}΂�R���394�
�^�fY3��^/���qV ���CZO�߃$����ya�3�:�ŕ&�v�=�~vo�)��l���{do�,Ro���o�+��MU�[_i�~ ��8��&�X2��z�lS��_w���O'���q��`[��n�L�!8��k)�ݡT�'��B3~�$��0>��>9��+��Z�q��$�����Y���QW�dY(���/�0��p��%�m �T\��̷� ��c�wE���Cq��ܦ=|F�Crn�͛���aetq�i�cI!��R�Bz��ا�^-����-��߲��$��S��ƃc;q��B�aѡ?��������DM���13����M�c��V�v��o��w�:��qF+�=v5����*� �kҺ� ����@C|��!����t{�Lx�r��e�eN|	'!��P>Ҡ�����G�G��Ĭ���K�S��U�Gm [�i��H8�4 ��25��$�����%��z�dP��*(����=�VI�!,j�3�x��D�_A9���ou��E��#����[�Lw����=ו�aA�o���*�U߸��'|��u�Qe�?s� X�9=����~n.p���b*��Z*��SROkb�HoI*�o58i�;v��!���׎��j�zǅH�`�9+��,�I�:�`�̖�ҋ	#8!5ɩ!���Y���
f�<Eʲ��MT=��$�1�xM9���U�������9�����;ڟ�y��l�h�ݫ�-{}].d2��Rf?�5{��;������d %�U�8�D]N�£^�Ӵ���p���EGc����1G��<S�V�릜�ȁ����\������������V�]���l%�b�/A�K��*C�\�!(T	�qcfj�ՙ^*�1*c�p)����f�y�*�eE���^���8��5���Ԍ �Z�X�#!��n��n�G�Yׯ����Pd�>�����9X/�J�4r�D�Qk>���������7?A�M	��V�H�p�2���S��0��K5��.�>��[+�=��6&zJ����ﻑj���>*C{q�($ɟ<�4�Z��5ɡ��r�mW�+����|U��idb�_��h�����ʗ�~֣�ɫ#�J��X@7�Qͼ�o�1U��(`qg"���1V[�K�(���<`�	J��(~ �æn�֭���n�	"�80�Z`������,Q��AoT���'���FP�`��[W���2#zq��iq+�L����*�\�I4�|�'+e�O�z8�#-ʻ���gk�U� �D!oW��$�p�]�4�������������^����<����t]���\,{	U��c�7�rTm7�Ꞇffex%p%':Uj)�aĖJ�-'$�90�]�1�˕��&鞑uw���Y�uk�K~c��-<�&h���B|֌lu>����F�8�"XU���� �C�͟B����8J0��B�4�d��Q���r����#�WM�"
[()�?IƲN��1c7-��h�uU&t��s��x�y7z��s;C�
��:�?���g<L�9h]*�B"�{\%�m�N2�����[Ju�S#F��pd��'Y�{Xd<�0q��֯�V9�p�Y��h����$�>�;ː���A$I��������;�d��Mx��8���|�~4�7r����Z��C`i��m���v�S�Fi�/��au�_F�.Q����`��W��+�*� �
���Pc�	9h�k�i���Puo��S��mLBwλC�XM�֭rɭӭ����ra��|�V����3�r�Jzx_ ��� +�>3�LB`�K4�Ui�L�XlxVHYEB    fa00    18801���HmIY�|�E=�g�C��cX�
��X8&~�����w�g@�%:�T$,x<.�QFrMv$�4?>���VYo:���K�)6�DI����$��+p��՝��xj;�� �:Cڹ(q�S�]��< W�����r���f�Rk黲h�&z�Ϻˀ����Zw����E_�ws����G���$����Y��I�ڱ�P���x&��g0���� \2D7#�ū�](�D���|�U�Yqг�ڇ�>��j%*��G�tۮE�hc� -l��0nՐ�`{#���6m_:��Psq�p�ǒ����fSZ����n��ڃ��1.KDo��^��7�-�0�TߓGM&�]�Ƣ2Ϋ{�۔��p�[Ǿ:ld�-��h�U��J�u%�k�y�t��$��LIe8���[ R����������?v[��<LM����Ͼ^��@K��<�BXA$�&?g��[Q��!�u�R������Ԅ'���.K ���y�X�h�5[92u�2=���A��_��|�@W�/��86���	��2��r���y��&{�b�iB��-i^Z��li>ޢ�����9��I������g/$�τ'xV�M����.L��C�1�2��b��o����d;�adj���#���'D�-��#�j�Ȣ�����v��P���:�}ق�����6�#���3��sӭ8��L������g�jJı§�#�-�ej�A��S�r,�o]a ��Hi_�\g��݁Oxb�t��Rv�MO1�,?����ɜf�)���|��I��x�"�\e������+����T����Am-��#'+�}��I�}p6�T�{��%о��}�g�	}�3;|4�8o=#׋cb�g���ۻWH�}^�R3���-2�<�(�<���y�f5rcP�m���<-Pf�DF~�N(�e�8���0�w���YuH��	2�2���Hޫ��2�}W2=Hl�b�Nw;�4=��T��X���ڸ�v�j�X����/yZ���z
}[��\��O?�>,�'��znx�߂+-��b8�W�,��d��b��Z�_=4�������z�,U@po$��f[ �������N�ǒ>%d� &���{���}X��p=��U� �y{�gU�I�ސ�k�)�]���iA�N��	ŗ.%{��PB����בU�-��;C��zD���X� ���������s�!j�ԡ���>�F����-�hp�����C1�Xw���8L��!t�T������������.��?��]K�~��K�B�3���#mQ�O6x7�y����G0����W��h�7�BZ��҅��_�z�"�3g�a�;�+���b0"�'��Ϝ5Wf׿C���D��W��k<�g�İɷD�k/�l%�jƴ�/��]�{�����b%c�ٙI����ͅ���.6�f�N�Y،/K�~r3��h#����Ə��Q@��]QA����Lzfl���O7d���[b_T�;�}�������?(TrɄ����B���<���+��	J�>����GS�v��q���6/��~C��j�ngq��̫����'M�W�ew��:\k��Q�v�52�c��K5��70�8Z�x�.s�����z3m驡�XH �C�h�	Q*��z������eΙ�䐺$vT��4�& %�A�#G 3M����L�]<��d<S�4��y��W싹�2Ӣ�\��?�I�_���'�Q�b�S�rt#X9�B��ȁ�>�}�tڵ����Ӌ��C��I^T�r�V@i�^�w� zxE8Ew��sc߬�s�P&g�`C���'�(������F�*�3,08	򈚷_3�4l/��HG�Q��W��jXhB�#��MF��UB{?�g��&i�p�o�_o�pnS,X�P=S���*С<�����5���x��F��֡e��q26��"d�b�P��;��.�6�#�O�R=�G��-�B��$�T�9���ЉN���� y�a��\�8���<��gc�������F�1 �~Q��A�}�$�^qҎ�v������ߵ7��e�u>�ꃍ��#�9P.�eg��vQ\��3GTvs&��z9F��;UÏ�h�Fˎ����G��<$��;w_jr~m�Y������l`U��/֐��=�%޻�Q�@�g帽,?���ww�ZUM�E.��h�Miiz������b�w/2�ͮ
�]��f6���z���',���e}�Pw�ԫ]�N�闳SךC��]�2�G+��PL  ��X���
ENɂާ"�\��D���7�����K�CR�V�H���9)�eĤ..<jde�J����t��J�5��h�Հ?-�������#�7� �^�RBg��8"�U<KՐXRƍH���8��q�w���px���V}�r��q�M_�ø���� ��~
c_������`g*�����H��*�62a�0d/��}-�X� Oɼ��C�T�v�0A�Ϲ�J����͍�A�Q����d&|¯\R�o�k��<46�m	�msX�ű��^�v�����-\����N�/�Xd��`#.J��2਻xg��#���ݱ�tR����(qMB�|'V}��D��fȼ4�)�O2�6٨�|/vsr!��c������i���qԎ`���t�������N[�o=��v�7t��bJ9Pb���(em�5���\��gd$�j����_s�X���(1��x�~N�8VK���7�z�M���
G��G+ǝ��q[��E���N��yIٌ0�k��q%�-�$���G�{z��񀸹��]CD�"�U��TEÑzy�9#�FL���i+UuW��"��󫆴�ğs:�+��]���w.ג�bN��[��{OF�j��G�ގ��Kz��B�+V =��I ��ͮQ�|d��+~T	�L7�Zf�%#��6�4���A*�<8�|�z|cyw
�X=��e��Xg��*���+�;;���,�uҏ���S�&��K�����ڎ-�`+���9w��1�Tj'	�e/d�+n�=�Cڗ�X"�0f97e��:C��+����Ӭ���c�3�%��h�QK�@�hժHk�y΍R�C�u�Ba��o�8%ބ��?}|��7>�O����>�|r-�	�j�k�����2Ⱥ/����CX{�'���)��:�:�N���I�&�oJ��ƽ���+�������7l��\�qz������sg\=�3
��i�9�>��Q��Bf�~�m�����O�_9'��#�k[��� ��ZeX+8�̱��iI����e��*���� ���=���5����X,f�n�P�o�t��*��8�*bh?sH,H��r��J��>G�� �{=�US�Z��-C��?j�{ӢkߏF/zZ���\K�G��)��iSBѠ�l���+<4�W0
)�4�ҍ��2��>}�⚫	�Bӟ�;Y;`�<����ؾF�kIF)��%�������䐾bV';�>F�����P'$� .���rd��u��2���>𧳐���Y�	�<O�������+pX��(�e�����p�� `4��%b`V�D'Ԇ��/.�eD�1����i�Ev��p�\�?��u����
��w�gt�w�����j��7�Ί*�P^h�Ľ0Y��/��d|�AЦ��v+�~��JX�"I9�^7�p29�=\��]�q����RJd��ͣ<��:<����V��|�rF���m��O:�e�i>�;ubXG�B����$�G�Ŝ�
s ��6�Gqn�_�]�\oH������NDL�Ts 2�֛�X�o��^�j��k;!�09����R��%��ڂ��%
���tM���
i��'�Nk�����͸	U���
u�w��8���"��k�]����{����ʏg:(�S���LYDi��F
��t��PZ� ����>� �~�5�c �����+a���a��,�+��W�'�\Pl��.�Ň:�n�Ҙ�����O�<*
>��T�T2c����I�<��Ee��'7�{����ҒN�Fb ��;�WJy�7����X�5�}���']!�o�f6��ܯX�5�2�c�P�U�E�q�^}�Q"���Ȇ]+�tǅ��4G�����������ʃ���M~��H2�!E2u"��bSe4A��?jo^���Q��}�1�ʫ�*�yw��\�u��(Xa�r�en�%�\\�19����&�#��	K�[N�wE���/�("��z��DNW�ǶhY�yPT�-�k���6c���k�9����tBMlvί�}�g �ū#?
�)�#Ϫ
c-e���z��i"��%T����+�����(L C�"�5��9���G��V�6y��o���/KA��`�8F��9V]2�^�k��ݡ�;�^�`���'���f����R�����������$/�-��i6g����WP�#]�T{�/��S���E��Ƞ��Y��bh���;��e��_�J�A���X�Ba���~}n���2ۡK&a�Q����v=�-��_���+}��Ӓc��a�u���q�kw*���o��ҽ���$�,H� �5�a�@�ް5�Q'��c��j��I
@��>����X�{5�lځ<�{�[���R	g,�T���,�������9�WsI�1�~�s:=i�d���e�5�I�Ϙ��B +���x�z,��[{3�x���_�?���&��O���R��h9�/�䫝�i�ߕj�vU���r�1E�P�롱<�lW����e��J��5_Op�Ne�7�|�Z��,���%�v�p��z��)~$�9�ɃءP�4���(����2̵#��$�;��07���7߆ɉ��u>WUM�w�=�p6�;ך�ܔ
z�1�J{]WF��%5�W�_���❳�����3�kbI.�{��h��E�L��8z�Yϊ�ݵ�|�t�[�p��		"�=��T�܊͙70�U��x�u����P�;�Yo}a��7�#	�.�B�ب��A��'����,��g;l�3G�aZ�h21�{�� MD_g(A+��Әn��f1b��������'��+�փ� �]j�4�FP(��lF�7�����%<�����'�6�k�"m�"��洩�Aa�K��mhs"��D�4����R�3��b����_����*qM��n���X'���j{�>�$j�OM��T�'��v��1 �w������� W��Y�V�l�A	�믶���lE��L{.���e(����>d��!�	���s���E/�" �{Z���?�	0m�F�.�{D��%�T^�ϖ��Oh�)�|{S偱!$dC�(�D@"��Հi�};����a�t�x�O��J�h������z�=��5�:B�7=Ց¨��I	�:��������5����εvm�*cTb�u[����;�^�@Xd2 t0�#,j]%r����Ư{҉ۏ�$鏑�|�s�=���r�7���Z�@�)�B�˽�F�n��!���v"�$ݚF�ڔģ�s���t�L�ўi��@����.i�(�ڞE��U�eZ�ߓ�2G߫Iך��NN�"���O&W����Pm��a�
M���bk�gg���_��}B�9&��9�jwW��|ێ��,��_ب��3
v�b�`���Kjٛ���~ �QH���k$&ݠZ`}'Ƣ��h�;�̗t����n�=�q[���^z�[]�'��~8��/�z�6����^t���m��d�d"���*|��3-9�+���3�`�G��<v?&c���N���=t�fv��r������H�M�u*SF���d��u���ڠ�Wel��eVՀ���4�i'}��Ad�!���Ը
SQ�1m&
l%�N��c�S�.�Ǔ��x>�����'(5N[3�%x�F*�?3R��(��|�WF[�=�z����W
��z�ki�6�n� �i)T��YJj���^'d �o�"޾D�:w��U�W�daB�<.2�:�L����H�1��@J��%�T{:�9u�0[�v*�@ڊ�q��N�T}N�G�_޺��E��%�{��:�q��v�S��[S�9Y�K���J�}h�IBʘxۏB�u��٪uV���fy**��\�[j��!�ƞ8�ߗ��j�aP�T%�0x���XlxVHYEB    fa00    1910J ^J��n]�=Ф}�/Noo�i�	��D$ޣï���pV`ތ�Q�T9�'8��F���̱����hZ�1jl<��+!l�q�Jirƻр�|���M�V�T8�<젖#� ��'r�X�mL�'��0_�E��υ�8¹��՛���8�|ʷ��(��DR��P+O{�����3��"�i�1YE�� ١CuP�O���%�XH���^^�A�5���/ua���rB, ��7
�E�l�?�za�[w�J�@(��2��_a�H�cJ�7I>}�(�	�~Zd�'��5�K����y+�gy�����J~,�r�ɴ�������U��^�����
�t�rdu�$�x��:~����*K�f5%Pc�nsYG�i7�����YS�.�8{%�e8W��.!�5u��q�J��������Ã.���M`�u�W�s����&d�:M�֯(����C�����lH�0���KY!o�������Fj���
�?�<��t�1{�:u����^���u���Um���� G���:O�Č	��~�4�#���׍�f��yF���\�B�+	2o+I�ֶS��V�p����6"d����gD�.�	0/d��]��-8r�$>��j���z�nl�+�\.���%y.�'�lT�f|��1��G��������EQՇJ�#��ߵ#;"W��[� )���wu����ơ��zdW�8�A�%�S��;��2Y3%���8!Gz����@c�#.����8�]M�q��c��GҞ�T��/�E���!c��͎�,��Q��$���EX@���0)i��C�F�JG�WH��n�++�C��@FdwLg%�D0����2C1���������/3�`&r��<Ǽ�T��9�/9S�Y��K�,���D�AZ�M�]P�f�]Z�Q��&�u=�����w,czz�S�.H�=v�v��V��)|I��8��� O�(K�<�׍u����,_TG!B�����ߑ�V�e�|]e�@�O����$��F�hw.Y�?
�!BH���g�A��]{���ܵaìk��� -ίR��g�$~;���ɟE~5��L��w,_K�T�d)���i��K����z ���ՇZx����q[�*��ݼ����ֿ�BK-�ڔ��:�_�q�����b���d�KN�nǧ�0B�C̿�GF��������(�=)�O��k���d�X�øʠsI�)�*I�����T��j�z��2˶�mk��
&�·D)�2zw�J��K�q���Ζ�^�~�ِ*�T��b"�\22��vXA�ΐ=ǁ ���<)�;�6ܑyG!�|��?���X� �>��ܴ-�z)��!���g���3ߢ�C9�E�'�/im̳К������(2,� �.�Hͅ���%�&��E;��$�c�2�W���=q�]w\ �g�tם��A��C��l JG2�	�Ɇ����bę���^3e�e�i��-����I�oIx��l���L���{(Ė	J�Nyk�(|��p���P����m��S,��[��a���[	H��6v���k^�ކ�'٧6�k 6��Ô��Hf�B�3j�Jj��&v"���j[��dn�[6�q>�����![�C �-l+�?�j�PR�LO5�|Ӽ�ѣ~��G���;�TWn׵q]�e�2�	_@�������Y\nŶn��4Ƒ|��Q������`�]�Dȥ٩W�v(S�G�2�6���q���$C�*��P�GVg�,S��B1b�{f&�r��he�^����Zd����gF�c�!i���Ð����k�0���57��r�����"�C�s�Ӏ�����2/J�֚�S���Б2����$}n|B
��/P��2�$o���{���jAh8?���V�i���,�0�؈��y]�% �
H2y�HK���
�q�J7[Yӿ=�`�R�(�&y��?��aHO�q�1=L
 ��q��g�*�ћ$ƙ�c㏣���^�P�/m�&8㵻3�n},��J��H���@�*�	s��]��UBQ�j�pv���:���Dp�=2!A��"�B����i}�$m�X�D�4��(�3�fT��HCsLI�qe�V��FW�1w����w%`&D�Ӗ=�&H�-�����L@T\�➋eu���/��tctތ�\���u���&�\��/��v��2\�7I��h�B���v�@���y}`��p��r���Ϙ�`��A��9M���f+���	�i}���_����Ȫ���v�J\s��zL%&�hE��vW���Yw@M�Ҵ% ����)�_�۠]q�+-C���l�jFl��U󆈤f��-0�����#�A����wîd8��0ٌ��������w[1��K����aY�QK�������ʥG4P$L~/ў6 ?�-h���� ��#+�fҰ$W� �*z�Ҡ�J�*)��Ś��ig�l�;V*���+�O��g�Q�j7�ҕ����a}��x�#v���`_�v���/�$5�S���"�6R~�_�����툔�a�:|�5Wap�z1��7�D��F(���>w_�*�;�������8�f���U�S����M���ʯO�P",�5iq8�g����>�O�8�-��-7%�дU�*�mT�����b�ԡ��c�;_�;���.�#5�?�;KM56�����M��2u
���G�Ƚg"ͱ󌏰�-d)\R���!�}�&;�$Z�:��T�?#�{���é�1laT�F����gi�@��O;�� ?�N��f��Y��j$h��!u������~�B��P��=d�F���'��f��dr�gAP�+�u��{Q�5��f�À֨>J�j�"h� �֛�ہ���t��I���,��j��)�Żry:�8�8�1s��U���1OM �HI�r`�>��x$J⾍W}:�7,K0)-B�*y�e
[)�XD+���;�K�X�Q�x1T��鿚�+}3���i�)xb)nڥ�M)��V5;���CaS2�Hg&$�o�$���0Fx����U*�/�\������\�������G��_jv�]��������VR����������,r�|�g����'�pmg�c�<х�MZ�6hȫzs�g*A���@?7���H(�g[��X�)�j~�WJ���/�X:��GgI� �wg�B13�� G���a~�}i� ����Kp"��O��y7�MS#s0݁�\�H�"�t���Y�9J����$����2�L)�d�1izT�?�}�X=�J����ȑ����Id��C"�{���mV��RF�1�O��=٘���f!��J�\�,��.�W��6G�rCD��~�����6o&��}�v���!Jg��v�L�}�)�6R��G�	��l���F�K�	!��3��+�!W�Û���������6�o=9� ry����X�<�P`�UZ,�u7I�����#9g�3	
����PU�T�*O���'����!! �|���Ŋdc(�9�9LQ�ڕ.���8��[�{ؼ��ߝ*������y�Sɴ$5�cc�*n$�H��"]�t�V2F�+HIˉ��w���K�kD8swt9w]��S�Y�k�$S�sI#Be�yo�)GBD%��fT����8�Slx<�Aˑ���`��1q����Uy j^:� OZv %$ ������^A��h׫)�jN9��õʗw���pAB㻃O�jR'^:����3�A��{(Q���б]�����䛛f� �( ڀR/�8����Y�F�0
��P姮ئÚ9M��k���C:�Qс���!��݈�:�5C8�Ia�Pv����1T/��ۛ��n\Չ՟��P�+�R~0�;f���/Z
t<t��m��F�'���D ���Х�#V(; ���$+���hc؛0���k�P�Y?�� 0�5�m��0*��r��P@{�,6I^0YX�uʟI_�������K��u�&#<��
mY�bs&d��'��*Ц�GkY��.���k&3��|�=Y9��	mg���A%����z��Ϳ`�`M�������$Xp�����P<b9�����(��uR.�����qMA��:mc��\�8��aG�%T��c�g��X�Q F�/��d2�N��k�����	�7w=0����J#:�������ê�׌��)�{3*͙;��w��Rh8ͭ`�J��oH$�!-.���x�0q�5y6�����M��2
.�ݣ�A�W�)Z��(�&�U���q�V.2�� ]��M
����6{Wzo��LL^ạX�]ռ�s5a��(ܕe1����CQ�9L�{_��k't�L��d�D�y�u��\Fң��e�+���<������ɠ�Z��"� �t8UxK����&��}��ͩ����m��مl tK�	�l�
�8J��ɱ	�MC����"�
s"����$��1/sG����(0�����U'¹	ē*�#�.2��͊�;<�."�v�7+J�z�A�:���cH1��8\�o٤��ښ(қ4c�/��������Yh�͒�T9�E� +d� ^�i�Ps��\�K^��/�K�n��?��K�6I�[��w'�wg�A]�S�&���^�.2v3��#,T�z�.�U��N�{UP��
�����g����/,ʴ�cz�*�n��҃=e�7�m��\( ��h�.8�
�;�j����^��7�^�O����c(b.eL] �Y�g����:�;r���=��o A���O��i�_�W Q�m�E%�W����Z�r�������٧U���`�}���mee�ޝz="C"���J�q�Q��jṥ���ƊV�,m�e/(;S�[XW=̜V@��A�|B$�[3SrĨ��_A� &/?'�.ӣ�i��5h�-WP<�,�
S�5�F����:�����ηɩ����oHm�K�<?�����y*�a����(}S��./�ۛ�=�٩W�I~ǡ�OM�A/���~��P9`:6K�"y63��-�*�AD��޼�vIIp���?I����o�H�עN�H3��_i�xE�@c<��d�jl�Aq� Q��Q-@`=F��9Z���������|k �mz��� �^���6�V�r.��F�o���@Ԛ�(!��*$ �^�[�7�bxʋ'���С����������d��~T
����zj�Bq���	H9D������q��m��^��#�xJ��D�sI&N�����9��Mmu�Z<��$Nj��Ȯ�n
e~a%MG�@S�r�
u�d�i�����¢��UO,�^�s�f�HL|l��l��Y���#��9���l�U�At ܖ�UU�"e6]�Ǚ>9�duPk��D�z�c�uT���<���C3��|K6��	���o��O��k�K��
f��/���Q;��8�b����������}�Z�(hy^��78J�欑�{�����czXX�qk ��D<�g�;k�X�f��#Kk	���JH?�������\ 4Մ�l"��ƭ>�9��W�&	�Hh'/_GW�ze���=���%�����2���X�@�hTO�
��CmQ}#[���ٴG�\��BUF�7`����2�e�'�l�Op�%�Ƙ+�@>��dKR"��\�ڴ���?C��y	�c��l~��g� ��Q�qҢM�y;:��lY�W:^��+���^����/�3h���|�ՅI��41i�9��#���`�s��(`:��v�%�?!T/���s�v���N��һ��V���2�<�5�\�L�Z�����=��	�ϸB�)��մD� ��5�獄0?D�ZL�$?���t)	��'4놴E���N��J�M;云�Q�T.��5$5<m�;���W|.��'�{A��Х�8�+����I�W�x��fR�T>p�}���!��W���|l���mrI?�<m����Pb�X�I��L��*�D��3�m�~b��!whB����6��D�x�]9��AxKs�KQ SùG5d���jz�<�1�7�6�	�u��|�ϡ[�o�z�+r�x]�"m���ߜz���9�W`"z��`V��GƂ��eiU�����.�rM��E�����΢��:	�k���R2���h�t.]H&�/ϡ�o�9�J9�_��T��PV�|J~���c�Y����H�9R�9p��Xr#�pM�8��@D�O��p��.���=�%�@CkB?-)ȅT}3u��7O�:�:�rK�q���W�t=�ɼo���c��U]S.��!P��%�%��Cf��4�H%r0>Zl�4,޷�Q���G��\ۼ"/6����X+�{�85w�Eg�@�M�QD����\)����XlxVHYEB    fa00    10e0S��K���FM�3�����)lw�^�6k2��0�����b��I��hB#B|��!�/g������t���>}�$|��Kr��E_x�u�?�Fw�mZkAl�c�dU�B59��H-_BpA����#�+�x�Y�����Nߘ6�]��7�@ړ�fPX#uFJ�������yܳa16�*0�II��=+���<���9�\�v�|�|.��D�<H<�d3��"�+�*�}-��}ܛf`g��l�W�����|a���������5��-8WU�&��V�"4@P�1*�ɜ���kH�:���	���#�����9#�Fws�X�kQ��6��Cʪ)�ɶ#�d;�֌�FY4�KQn��9�j�|J�5����[f9�b%��.~<f�bx9{�P��Da������:���b�*��|�wD+�ׄ[�9��/78F{]{KK2�fn���	N��y|�^O��LK,��ƪÑU�5V�&��k.��V���%u9��A\���}���֛�����ԨT7[��A��L����{<�C�)�`t鳄��/�(w@,����X�>�O�WH��χ�������yf����c��=�΄N~+��j/E���p�ዤ�qw����9i���|�M�E�˕3�OQȿ!���nT���AA�n�Ql��$�q��]��e�S�`�������	��P�O��싽i���_=�f�p�$�k#Pu�����s^58+ty�4��I����H����۰�i�A�Ξb���U�U6r#�X0m���vtP���
�p?��)��HA�f<p��Hf��f��o?x��(G�GP9V�V���G�X;ՐM�+��&�mXpK���C9��\�8����^<�ѯ�P�|9q��0�����M�ׄD�X���.�O���<�d_�gͫ@
v�^'��};�2�Ӣ��ٟ3xծ��w��ԷW)h���#7��3�ݔ���"c��l��vm N3N8�Q�
Ś��b�8f<w�I@�+�B��xm� �3r�;|�S��]�S���O#N'Cȹ��qW����3�K��$,Uz$4[�3��m��V��,�Uv� /ٟ�����=E��~�/3ҋ���$�Q� �78��������O���I��+ �؏����u�gb8 c�ݩ	�b� Ͱ��O�B���g��^2�Ë́7J�e�V��2���w�5W�l`_�	�[� 'RV7�X����i	�������H��Dt��݀�*���Ca����wk�c���n��l���HU׌�L�䮛�TJ\Z�H�|�����CH3�k���C'�>�wj�-.ɍ�7�d��ถ�E�%d��2��痙�/w��J�q0�.�a��b'V�++Dq�v��R�%�T����vՁ�b�m��3�4<�ICd��ڡ"��4��w�"�F�,P3@�f�r��/��O�H4�ċ�W*����c���7w{��=��Ц���m)��5���PQ�x0 g�<;��K�S��+�h��'>?��@�x���!�VRXu:O��i������Y�e*`�5W ����[ �%�&��@�=��5f���LI�:��i�:\�4�,ݶh<zx�@�)�5'���j��f�w��/ü�����
��ɸ&�z��^Mo��a��A�$�r��J�!�����{�*�{+�Z�@N���6���w��R,rЫ*.��ׯB3�?5��7#G�~	�Hl�����ύ��6�Fԟgԉ�;M���q3����4�� %���@�+(J"T�]_e���5�U
.�T��U.M8,8x{\��P/���Eb}{ޢ�M�fUd�;�a-j ]�ѵ~
˱!brH���V-O+CWŬ:�=��7`Ҷ%4����>��TZ�= uP�������>�־��L(�A����I���V��uZ���i�~_9@�sm>V��}��Hbh�h_�O��1�/A��[P[�W(xtU�Ӧϳ�������r��x=e�B�e��P�4���[����6�m`�	���tGM��+�l �be�M��edF�L��x8O�R4���gY����^�$��J�#��9B��'\�rIoW2!1�S�~(��fe0|�ĦZ�Kֹ�M��q�_k�g�� d#��5�
���V�`��ůe��m�F�;��C���^��є@P�y �N����7������O��k����u���zz�@����o�z\�[��R�%9�a��b@շN�+������A_�2r�f�%��A�=�� ��"��t<S,��/?�/[�Q���L�=?�:���QB��l�4��7�Yt����'A#���2���'���ʒѨ�i�G1�����m���w&��O��e��4�]ףʀ���,f���}�G_��J#� �:�Y>��W��+����]���L�H["<�p��.s&�Ҝ{5J�lpx�L�듟� \:@��f��?2�%5u�[�����M%a~��݇Mf�8Yrd��M��=hEwU�(o��F�yc��N�b��z��p�5 ˵Ȭ��n֘�"^H0�z� o��g3q4%����?���G��m�(M�A.ܯ�{�az ɸ��t�HL֟ˏ��9|���:��1�ܫ�g q�ۄ�[.�97	�4�l�+��t�Rk�M�&16���\�x�Ә���@���Nq�����j�)*oe�E2��������p�P��{���O�_ �hk*���?����C���t����	1!�E�(�$.�|"�۶��,ƙ�GG}�G:�n��.:mJ1�
���H�]%�������3}���@����;0���r�?ѮCAVy.S�X0f��n%فw�9�J�u��O���b?�� D!�j���:���:u��y3!W9�T��%�Q��G	b�Rcc���ٺʹ�2�S��g��E��"Gq�*�T��u��L��@�j��Y����$z:k���w؅�� ��T(�;��J�
ܵ��YMt�^^vx8�hnhB�
h�y��G�J������׽9Ɖ>����`�@��M2�ۄ.��6I۵�8�z:����_���'\ ���.��-��u�AHo�$�4ʽ�	��>��R͡�p��"'踠�'mc򺒲_��Ꝇ0DM=,}�Z���ːM� �K���*J�zvT7uxjC��=�'��ƛ����t{E�%�1���b�f��@���8
U�����3堩{��~�k/�.���c"��,��a|�0R;��C�P"^!��i�q!� h��9p�oJau��3&5��%�K�tUw�Yy��0KV�=׉{�w�K0S��Cݺ-�8'uF�L��qU��(+�+�򥃿�ÆϬ�C��W\���,G|��R���P�~<�
���~��
�q+u<_jh��*�F��0sw�G��߅�&X4k^�� <��Q᧢rd�A�
�IPN�7�Ls)���t|�I�=�T�"���$&UvH�x�g􇧀�56�>$��d?�m�t,o4�H"
��,#�h81w�
 ���+�v�lH_g��Yʶz��|_uEI42>w����}���	C��z��:�s%)2��ٗ?u���-m�1�K�#�9N��D5�ZqR �Pi�hn��8��ܕ��=�"UaIZ��?��Nmvɖ���?P<iF-Ъ�nm�,Po9����#{O�v���X0޹9dWĻ�8�{m�hP=�ԯ����e�yjr�BL����mz?��u>,wxf�\6#�uY�S2��Gȯ/�B^\��EwS�m4:'�l t7�ly�T�uQꧤٱ�1,�~�,��j%�%����(x<���h��R�Y�6@�v�	�h �ٲ �� �+"Zd����u(���ͅ���O%�I��t)L$0mCO�:��Ν����H������$�Ά}38h�2�c�p�.1��ć~鯋b9X�vk����b�������ޝ�.����[2��'��G��S.Å�P��e���i��7N���Қ OlE�Z@�M'TI����
��,��f�:�c�=���������Y�S\iL�}��rMY|y�x� �>��}�-&|ڹ��/����̌�a$��ɧ��S��#��L9��$�4 Q���UR�ڞ��R�[��+�i���	3�.���B�f����nXx���z�R]8��^)�"�%�t�_�&�'-	�d��dş�����~HI����q���͝!�Z�pZ9�[�l��'�bf1[���0Qq��Jln�u�F�h0��cy���Ec����+���_b3�螄�Ƽ��� ��I� �XlxVHYEB    fa00    1860��y����Ɛ_���^:�[�ԛ�>Z��E�kG��-�Ɛ��47�2�ܽ���.�
��3O�N����f	�y,;�XE��8}@W����p?[`�YO����I��ΰ6�<^�q�狜d����y3�5�P�f6�W�KmzR���u�M�Jp@}�I�^U";�
�B�l�d����#9�������أ�<�y�k�2F�.�Z�c�(��Y��F!z�~�vh������a/S�u	o�G�zԍs"*��oit���[R��H*�l9$��b���	Lu�����%�bj
���1�d
umk忂 Djp����퐔�l-�J����4���js�)D��݁��5�����y�x:%�:�خ��ew&��D�7˷b�;Gi�.B#�(,,�T*� �w����a��<%���y"� Z;�q!��G����:m���	��8�KٝAG9��D%Q��2D�[b5���ﲘ^��*��S��]����'�����9���
��3��g*v��DM+��L�}�'l�z�5ح�@~5�9	<�a�P?]I����5�D���eZ]�w���5I�t�5��o��t����s�mw60]Y��Dv`Cu���t#	�8%%���QV�xpX�@,��(��'L���J��CE�T�Y��n�Z������t�}q�]ˍ%B)a����v"?ɶM�L]��N��8���<�~�4ߟ��4���|5a�)�2����<K��8�lM8#�j�a�έ�
 ��7N�Ȟ��r�%�S����R
.e�T� ���D �"6Ef"�^���QЅu�	o��Qx`���8^5�p���>!lK����g�x��0j��`dC1�����4�f�&x%��	|K�!͈�z�4>��i]VM:�[�i��s�A$�ՇӤi��/*��E,���V���v��b�z�u>�Չ�������b��5����A�[WͨKTO�u�������lΘ��.H]�ڢ�Ӈ��x�Y���4�N}U��r�a����b��G���I�I����Jn��C`d�C�<�Ͳ�
�����G��}�.�%� c��b��Ny�ަC91�����1�ȭW�@�k���
��߈��W|;
W�x�Z��c�b�u!p�}I��O�^|i�E�j;Eu�̋U��Tt0>���p�c�[	��ݒ�GQ��-a��Ő�_��e�=!�/Q.��kk��M<;���ctX�y;|�"8Ity^<�}��n����p�X�{j�����/�?J���_�By��l2�=�#I
p�Ж__d��[�L���?���=���&
s������X�ES����	�wO�]1������ T�j��J�b ���X����ex�s=GxM1�b	����~�`�
)�'NnZ�W���9�������Qi��p�tu�H~�[QA"�N��� �UX<���o�$�,I�Ns�o	7�t&I��� �0J �Q��b���hpkZ큐�U:�.'0x���-x&e�n��#�}�6$��I��<�\>����nQ��#W,�u:�-nvsl���M:�N�nC�{eU[��5Gk�}D'Y�E�|��r�<S�Qo[or%���_ߦ^d��2��f(<L��U�%Q���]�C�; d������3W.�s����U�1k�F*���e��^�;
���~�5�3;|Um?6��5Nb@rm�
��f�����_2�1� �& tx^��=�S�����ENi$�ՠ�x�-1k3�I��I�T������&Ki`�\2�"�q�"B�F����������!3�
d7�}!����r] ��3�e4�d���\5[�.�i�L��C):����I~����M��'o^ٛ��?uWv�#�?�c�b�x�5��g���K��e�Ci��)`�g�B%��MN@��%���nh.���:W.�J?�u�Ԋ��@d�q���{�С��:��K}ݳy����Xg��.)�O�.=Ǖ�Z��\"fT%!g�@ ���	���8j��qd�!C5 У��7��@�Z����#t�f��Ө�Oh���:.|CV�J7���HQ���!7�P+&N�y|�hGr�ljC�0�w��c߹v}R%Z���t fpt1g��ah���a������J���]��U�lL����X���|2<d�h��g��_�'�d����޽Nc��A�ߢ6B�6j�ͱ�it�;1���2�B���F�� �c�+��~kc�C��Iʹ>Ѓ��f��V�hv���� WOn�f<��rQ:� ����-3s��^�	������Q���іAՃg�� W������)V'���[ĕɎB�L�.�.d�"y�>����<`�eo����]%;9��f��='�{���n�i�p�l����H?L�1����К�"�`�� �4l$�y�
��1W ����ݦqu��7:4p�&��ytJ��_J}Ij�F;ư[<q�&<��4A�e�DdU)%��2�<~5���˞�z����q�1[F�$�L�pa�c���pE4�e#�>o��L���T7�5q�WO=��y�)���0r��_:�����$��3|c��M	(>�y���\���ɏ9��Eq�mlC��õ! ���ҘӴ���&���<�1N }�G�7�J��H��`?L��ɛW���z�.?y�nC����Kv1r���<X}�S�r8|5���r�F�P6�a7~9�rl�5vIA�5.�(��08�R,��w`�~f�����Q���G��5}@�U�&o>� ��q�l��ɲw\�V���B�P���J�&���f.B�A���t���pX���S�6�� '��,�C
�YAtV(��w&��"�^�&2䄮s�$�阜g���E�õnqᠽ�k�CY��-q-3�DUZ~9��?%���'�g$"z0�^�o'��$l�K}Ĳ��yYt�������˪߭s���@�t�z 	�!�Ұ�og����E+��k�1�M@S��\��US;R�?	ݖ�����|dX?��~�s�JKo����M�Q�Vs����^����T�g_X2�r���ଭ�����5��Tm�?��`�U[�w�����,���;��Em.�p0r��3�{<��z���ĳa��I�[
����y�u�w����ћ�7�`=f�1�Sx������0iw���� ��
U��s}���W��^��4�I7	&��|�_#�h<������cɔ�ƞ��ӼEOK��.W�-C����l+:}z�=���
��C}�C��R��]Q5��5k����N�Q.�4K{�aL//�_�s]�Y�Vr榯�4Y�A�q�&)s0k%~v!�g������X���^8�����ndc�#����Lz�����l2 ������py`Nq���,ě�G�	U�`����7Di{����FAh���kM���
�����/��q�4��c9E�g���� ^r�D��v�)��{�ňM����L�&�`����9&s�u'�������zuoT$��Sܶ՘�V��+-��U�"�`FB�N2�ߏ�@<��oQ.��J���1������O�)�������|� E>D��Ig\Ě!4b�]�����~?��0ʥ����i���i�7��(Y�i]����-�.�[��������M��^�~@��<��fʜ槪�Bd(|�fN���-�����U_��b�+�&&��+�^���2ԑ�fGӼU<LyN�h\?)�T�+0V�xH�2uBtX^���Xk�x�>�@n�p��>��TI{d>EU%�
#D����޿�ъ����JWT��l�g����M�C�K� �0�u~75�\q�ٿc3�}<YyB3������<t.OY$�b=�G�SA\;(�Q^>��?�������˓nuE]��8J_���&�* l��yu���~y�'���Z��}�v$ǻ�$��X���<حy�k�p��{h������N��hRF��%�eːF���_��L���M�p��Rs��!�yM�})O�@3��H����P����m���]R="^\T"�H�gn�Y����|Gb�c�$�!t�?��"�ʍ6���3z������#��j�D��i.���r�B3����g�$	�1C��@�h9*Ŕ*yqg��_��pǩ�r*��N�0�5�\}d�^Ұ�Gl]؆�V���2"���1��f�oė&�y���RV�ɲ6��/u����8B)���V�����ZW6�npz��ф<%��\ó�&�R���W捖�"�rѳs�vn��X�+�ft�;n
i��]Ԯ���ķ�l����9-����-�%�F=��w�-�{�;�.PZ>�ʹ�Y$���'I��%ߧ��燡W�$�\K��b�r�w�.��,<��9bV���#��J�U:b���]��8�,�;�k�ߜ��KR�c:Ό8r��l%�̿G�o�bޞE;���s�VDa��,�֬�"�5�G�c|���'�H.���� �]�a�|{���x'ks(4:y��u���1�K϶�}&����۾pO�۔���X�z$�f�5h�i�'	,�J��x����@�z\��)����z�ñ2�A�o�N����iaL_���!׵�q+����2m�uЮ\{*�y:����/r��!9��=�q���]U뀗�Dg�U?�N�Ik"�zڊGn���B,��E�Ǥ�x��@��*г*�зf�)8+�~�q�#�������Q���6�"���~�3'��c����9��������ә���� ���A�T^��Mă9+���[,�+�a�r�
��3��q�W+���&�ݒ�����uo��N�T��� 3�#��,��!�C�����sY.����M>&���w�u`0�M��&/:�B��?PɈ^����jX� i��!�����l�+`��!}�G���?`�R��K�9M�K����d"�)փ0*��>��c+G�=A�v���I�p	�*i���"���,A���C�<����Oi���3щZ#�/���8^^�)�\�@2�[=n���f'8�1�h�4�_���B� t��z�n�{��ZJ>�N�'rB�.�4���P�7k�W�N���@!����HW�; ��|q�f����j[/�qP��#�)&�qN��n�+�c��'�L)�=tPA�$F�xd�Y������S?	�Ɍ`��:�{�.c0c2�9K�lu�F
6�KG�*����H�N���Y�Q�s�X�n��p����ܣ��5h c�u�jV5H�`�/A�@lk�I��j-���Ȭ�|b��f�knE5?˪�?��� F.?؝s�:��ub���fv�1����&.|B#8����V3���n�ǵ����'/k��0��"�*�A$��z����O�>�˻ǅ�$`������Pg�.m�n+Ee}���,�lc����pQɊ����
r�� f�L,�m1fA٭@�6�>ˀ����_�2j��97���� )N���.)�]�[��Vdx���i�P��(c@y�og�����w�"��b�Jq�?��i�@mi��~����y@��LJ�U�d��ퟟ�3��Np����4Y��i�_�w�g�4��.��
چ�B�����/�@��S<��=�:U���Z��p&��nr��\�{j��8��Q~�NH���8s虥<s�hu-��Y#L(bՓ�Ι����x8�/X#r����&n%��㭁 �V�|���l4�}�$�1�fV�Z���䆣�^T<0���df�5R_�(ÖD��5����Ϥ��f��"�q�]�[6D�J,ۃ9B~5�Vz�����Skԗ,93L4��^K��I	��楚�#ЭzQ��xt-Ma��(9!����BW�u�~:rWf�Gr�~�b�7җ�=}�ʑ���)�ˏ�e����ʩ�H�^�����w�C�+��t&��!�}#*B�D�PD%C}�f��M׾�@���O0C���9汑x�Qi��^؞t֑��,�@�~+��D�Gv6���~�5�ؐ8aA�;JD��%=<�.w�C��L��+�v<	Ɉ����v�>Fd��kȭ#^z��t#_6G1P���� ���~,�dK��MN�~|t��Ke�yFa�i�M��?�XlxVHYEB    fa00    1720����l�#?ʑ�Dh�90iZ�iid;��f�F�O��r�!XA�n��H)���C��ЋKNț��S�$^��u��*c�N>�R�E'm���F8+M�MU{�2�������6��p�1�����.	�Ow�v�݂}������������3���'U�ǋ��C��m�Q~�a�l�����0{Dd/�>	���( Z�it��6��Db"�d��踟V�bIl����퓼�RnPO@�U�ښ�K�2HD�MN|�m�?R��Q�wP�t)���cmK�M��	�_��96u�( z���=Ӛ�,>f���C
�eg�&���q�P�+X%�%������j-�ٜ�zޞ,hx`������nݼi�������lT'�B�"��DgTI�2�l���Y�����V��p!�87�ս+8Y"]���߃��<;)��AP����i�b�ܟuaM�a��j�+��77�����M��Î1}�h4�l����V�:4�J�	�H�>�Xo�oK�T����	�_E��7�]mm�TXe�N���_ޜ0�yLv���S��+��n3}�9J4E,�6=wp2�_�,�]�Œo}�O���!�n���BO� ��T�:h-��IH�%���ڼ`����� F"ӵ�)+;��j�P���4H��	������H�H2�F%�:�<%l�݆� ���(^r���`�l��l����a�dInX�\��Uk�p��c���A>,s�iy�4*���ʑq��/��p�it���Lg�m0���ɪ��wT��j"޳P�:�����i;xy�g�dEaqǻY��5 :��"�e��^�c�*�>�T�8�\��m�n0��� m��M�4�r��T�|����ӌo� �"`h���}FY\���[�<L�������3�+G~���G�Rz]N�xAj}ϑ6��N�9�m.f�)uwR�$�ȷY�r�ݖ*�G$�M.���%N�a]��d8j���AN�!W/h�d�Y�������C�B�En9^�_7rMpM�hI��}`X�����7���mDD_��4J��]d#s�kj�R��N�}=E��m2??Ax���=�+"\	�v��]un�̛�Y� Ҋ��tO����k��kQ�Bi��';E��	C���O�CL���3[��	"vr#%@��/�	�\���:���QJ3𻳤���:��ˆ�}�����Ҳ����R�TU�����H<A#�p��~�:"�1
�ɩ���q0ƻ�8Z��B�y;ʸ$�ʱ��͇Q���`�8�7ҷ��M Qi1r�E��ʾD�dGr?� �w���L~z~X��R�D4۲}�V�%���Eb���J���4�}�
Z0��l%`��~M�U�z4�8��k�__�{N��f���]v�^P�q�f�������5�0qN��a��q7ٕc0avrp]_pM3@ʥtb���T7���1�,�wX��2K���o1���j��F��\�I��k��<eG��I����W9��jt�%��c�i4��J�o��DUW�fur�ٗw8% �!�&�Q�R����&h1T0���z%ڎ��c��� \O�>�-���y�����-]y�@vл\w��2�t�X)Ƙ*�B��.R��2���>S������m�Nɥ����~l�rc�xOǉ�����fV� !�f��k
�N��:��.�.�jk��nF-�gQ�C�e(�����P�o#ΨZ�D�R)����死�T�Cs�/ޛ��WJݖ��&�Ε3鐀�*�#���p]�7G�3�V��;�,�]fK��I�$�V�v)�I{1��	uCpj�E������`T�%i���\���K����TӠ���Z&�~�Q�2���
Μ��:B��OH��
�5�My�"o�(�u|o[�O�73�ؒ�)�Z��J��i}�1n5K�F�O�"-p��^PI��:S<��8]Y����h��T�xO��O�}���Y��N�:��=mG�Bt�+��x��38�^OB/�9��ͅ}�_r����-|��d��/�}��s�Ll�:����J�M��	�)#����zD�92���E��4�痛>��Fs �e?Li ֌
.CO�{���;��l�k����V5�~g2���l�=�Ķѡu��S��Tf����ۄ� ��he�ǱS
�ZQ��:j����/vI�z���QK���������\������k��|��j�+�(�E}���E
�h[Ai�Hx�PQ��1 �׵���\���OGR����ٮ�@09A�P�
��@�/f��f�Q�6��Ԛ�l��w&���͜����d���v(g���E�A���@�4	;�����PG�GY��fM�󄬄�;,,�"w���"	�]ړ;�QԷ5���!a��Vf��_�n�5h�n{,�?,q��v��P���}��s��1�>���+e*�w�Dʧ�R����,Z���-$��)�1�P��RMeS2x�./��\ai��E!�TJ0�]�4 -q)�ܠZ�*�B�h� /̍����LQ�ۍ鹇ڢ�Eޖb�{���d��	��C}�KKDw���oz�L��>�a�C��v}�Z|6|�pC�c�ܩ��ӝ֣6�Z��}�ES��X	�h����50�HW�g`��x �%I=|�M/ɗ�a�_:x�vx�Q�O�o�kum�:���	x���y\��?��(������U�7������P�ڑD�p�A3D�^ʜ����)2Z�b�������F�O�c,HPi����r�bu�Fl:�8��l9�Jɀ�wѠ;���g�dz0>�����_���p�}~�e��z܉�7�
"�]|J9}i��<J���,�:�D5J��zF�a�/f���.�S(�S�%�!�g� J�6�N�/��II+�s���
�.�&��)e� ��g
�W�̠4�0{���֘�|X؏��u ��8f,kk���UA��R���ia�=X�C��<_���c�����
�JW�s7�!�⁝thM��/��4=8ƌ�{�~p8rm�A�������6�a�S�ڢčk6��W8�9)�i0BX�)}
ʄT��H�K�b,,�0o��٣v��͐��A��o����cM�D.A�Yo���UH��J�I_$�Z��e�ў~Ƥv��:��3̂L~��$��$ƾ8	���H>*�2�����s�3���,�t�1��mLj�K���Y���N1|���h�H�~�C5����L1���R�%�gVʡ����=����k%��'�(�c�J��vC�Dr��cH6FX����b����T���9����v��d�y ;v$�fx8�]8q3-��A}���b��B��G &'`�As[{6)K;ݞ����)�TꬹG�Vd�3\�/_W:7m:�o�CH0�����.QزnjT�� �#cX(�A���A�aɑ�Vgp�po��{��b#�N�']�K�/�d��� <~��
9�0��в7?�Ϯ~����3�z ;��ί3�A�g1l���n��2]��yl-�u�r�p�/Y~�Yc��-ΔwJ��(�Ù�[0���J8:�db2Jʓ(	�%�`��G���@ FrM^tː<T�>��?g��Ŏ��/+-�c��_bʣb{�p:$7��/i]�$�-%:_o�Y�.��i������ �N�nv^^t_�[�s�l���r��Fۡ�Puh\ZC���������&[����r<�QG��w�=(H֕Z�v4x~&�9И�)qv���׌��Z��>P@��|%��j
�}���`,
4���F��(ve�Wb;�5ΟC� ���?zpD_��@_�<��t�8�N�����'ӂ����k�O}����i�g<
F{�X)��^�۹6�gj� ɣ�����s�Y�n����3ʄ����D/�xm�����8:�Xq�0�2�Q�%̻�^v���l��JQaͺS"�׋`xA\S�Wo���G���rk��=��^�V��F4���\"+�g�2��$$H�:g���7��lE��
0�	�2���aM`�r�w ��p������NX�D�;!쓛�
E)��/����o�6F.Me�E�|���R�f�:��2p�n��r����B�V�F���1JD^t��������Q�G�ɖ��2�0c�6SEc��Ypi��a�����r7� �-�`����nVk��W�A�	h�J�8=������s��_�R��VyK��� �n��?���l�{h;��:Μ$bz%9����Q���NǠ+hꌑ����C���8���:��$��{7�1G�;U���՚���P{�%�f5߼`�$�Κ�O`����7��*�O��.�.3�!M��R���kr�pf�y�A9�x0���)�s[&J��Hù����޵�t�%41��Gi��O�In�7���)M��	���Y$+1��4*{-�<��B��^-�YRs��JW���f୰��"��A��$3�Y�>���k�hs˔N\�ľ�5��qt���'��%g\��)䒴�N�m$H�^�/�={}��Zʑ5"J��jJ���=oI<��c8Έ/�Ғ/�p%���ll+�Q�D��A%$���:�;���Yά��p;X'i�_��+qN��/+����&�\��~TW���N	D+j �V���Q��pǒ��9����Ji1zϽ��K˻6�K|bzX]�$��R�(��/���1c�t�#L6;4��يFaC�C�0�jDV��ظ�8�ʡѣ:�g���AGD�ٖ�?,E�����b������K���m�7�?��n�PȽ�>���D�J�_�(aM�&u�bC����Zyͥ���ܹ�"1כp��Rƌ�>�tL��%�X�7�jՙ�z���n%ď����T=܀B��ǍA�Da"i��yP�E��V����I��,�u��
q���0�\�ó�f��\�e˔�O7 ]R�]���C3��S
����cB�,���L!	0΁�����t�o�[í���9ѻ�2h؉Ωۊ"�l���Y#��쥐��a�����%�����%�EU&(���y��uך�n{�]n��_0ѤRm:� �Zq{������2o�xX�7@�fn��M�B+�,�7��*�����Q�gA�a�	�u����t�0Ed% t6"t������V�58P����5�����'���Z��kZQp��ά �!�M���Vj�p�X��t��N*�6ͣ�5�Ѱ-=����0�NK-��K�A�S�&�&d�C�+����W���s����U�fn
h�������ع���'��"���~#�'��ϸԹ2e(c�}Ǹ�O]�������"1*��0|����\��J>�k�C�NG�I�4�/��>���X�������1�#dI^�[ؘ�n���q�cר���C=�#V����w"L����6�����X(L�F��1b��c��d��9mT�62����*X|�VC�HX ���й��i����,LP���6Ew���<��=�t��[Jf���XQ@��$s�!��������va����l��/��ݠ8�4C���Q�J��y���#���%S)��Z�Y���T����,�.���-p�|���8�Ml��2�&<
�?*�jM��E3���F:�R{���~���Ш�t @��Y�)���f(a�����#�����M:�ﮯ��:��^aM0�$;;�	&�R|�_FV8�(�.]��s�Ś�r�/.F~�R(�u���$��,�J�Kx��M_�غ6��?����|c��K���.T��h����Y^�:B1�~�6�|�,����fu��U�f	"�$P�~�0�ip��h5�f ��b����҂W�'�XlxVHYEB    fa00    1500��� ��i_�:o�NV%[�A��(J����8�dρ�I������d�D�Ô��]xi;�pF���$�`�ג+��zl��Y����[�%F�ɹ�uVô/㦫fK��}�a�ar�D�5����Gۅ���2W��t >�^fBf%o�_��A�_�ۤ���'%n�\c�lo��!d^fä,����������Vh����(�B��o�ؐ+eYn&���z�Z^,��N�LIg�u��%�;^��o�U�J�	��lAL����)7*���'.0"�C2{`I���`Fb�v������Q"&?@�H"#��ˮo��L~j�
fN�sY���!�nI@��o�,mA�#�{ݓa�+�5���"\�Gê
Vc.'�ϲ-_�<�^��vy�j�GI��/�)����
��I5�����SM�0��H� LU��/	�B�2=�v���l1T��J=s�a�T'�$k��3f��G��S@|q��Oy���)��{[EI���J�a%�aJ��^Y'������;���|�0hI�Z�f���ۉ�	�Sw�o���_U,-�ǚ��"��{�Ā���9��8f�BQ܁s�T_Z�D6��ŀn��`+�#?K?B�O!�5ު��_\X��gN��M���?���������5�e�#tƾ����z�(���Q� �����_�Q�}�I���=�����k"�漭f<_��#֙����~`�'H��;���E�eG���!H��_�,[�]xp?�M�@H�R�����هjYb�����EK4��&_d� )��/�C�lPV�إov=1�8��:�|zTJ|��̜��d~	���l,���E��	��b&Ɔ�XU�@v琕2��D�1���:���qH�^5���_�6V��F�b��H���
�{�@9� � ~�7���L]�@�8!�k���P���Yq����|��`@%m��$x
����7�г���W���/�DyT�6�����N'����X�^����qې�7 �b�p�,j�Z�Z\����\�z{��䉼����"�fH�}��;�W@�����d��d�m�`�G��˂��x	lj</?g���CZ���i���ɾ�ʭ�M���z���d7`��uPD|��ۗ\��ڛ�;6�-����ܬ�*��_��ח��|�ly#21�rR��f�'L9HR��/�d�����ja��Wh-�I͉{F/��9	�̕Z�.:�:�BD�� �q;�bͪg%�_�x�����tgK�a��%�
�Ə:��)�|+|*y*e@��k���D�5�T����Uez�_~$�>�N�)ge\�q���`��Y�_���$f*���q��DAd��e�S{&�s۫X�����������6`7���d�U�;�4һR��"y��_=i0O��G�.�#�e�n-M,�FW��0�p�|,��H(��A����D�7�s2�'��gR���~p�rg�T¼�M^:���oU|~�V��?��ci��<NDo��L �k ����BZ5as�Z���r�k�*�;h.;Ģ	�1z@O~�o4�<�q��9q��Å1�ޚX�!�T����顲W�
������^g͒�}�����N��%	nt*�1���r��>d%m�*HF����=rɼc�qU�h�<�~��3��/y	�G���to^`^E-�X��:�>&	��w�� �83�Yz=�{}>��HP��f���BA��t�_}�"kz1���	 ;�b%B���/��/k�o\|
������&=�ݮ U$�\h��w������F�g� ݸ4�ň,<Ne	�=���y<A��z�MI�%c��ӿ���:��ّ�qZ��6�"��Z�>���BS�0U���V�	���@ט@���	Ie�w�U(�'�%��ɢ_�?s��D��g���21��P|X���a��׍<^-ƣ���\����b�����^���kކ��Ǉou��hw�6����� ���0_:��$s�H2<�~yvw%D
����%�T�~��ȴHMT���K�ݿ��H������t�o�UȮ�4��y�>�2���:i4�y�@F���cg��7�]������0��y-��XY��
8;q��[a��� �6�E��E�8�bN2*�U�wt�T�mh���?�أ��� �gL��ȦOP�6�[��l�)1�q���W�"]�A���<�e�����qk`ђC^֌89�m�YTFy��
Z�s��e9��燶�Y1�}C9Ϧ2�����GCo�}X��`	���&�a��i��q;MGD�7	?��B:/g�C��e�]$	���=��G`�gt�#q�����Z;7�I��G��l��+s�%�"�����A����]R��l�׈�f���f�l`a( ��&ߥ5�1@����w��7��_8��ِ'8s���R���R�V��J���Bp����F[�KTx��A�v�A��:8)�39`�}�	p�05�:�LP3��C�<��W�d<�e@���U`����ȝ"�?f��B�.�#���h��Ί�� ��G��]���4?��Y�y��W�=��d���d=R��훏�T���fK����!u�h�䈼Q�W��rq��j'���Lb���)��CTJ��\4v��}F�6�ixQ�D�������!�J�u$Z�)
��~�dt=�n\�57�P&��w�m�!����\}ףO���h(�Nmp�c ���%'ZY����X�p��E�%���l��%�!����#_4�)���-M]IEI=tU��N�qi��f��o$�42�D	J�G���B��e���eC�������ԉ��:p08aA+x�>I��������4G�5B��KT��J�֨0m����8^��V������_��R��M|���3t�+ �z0�ǧ�M"��.'u����i;\�m�����ålc⽱~�ᖊ�ʖg���h�:����2��DN)��.��Vi��4+��O�� �
7m�o���m ^s'��,���"��;��Ծ�V�i9Lk8tbR�'���i��+v���l�^沇ܻ��8���ÛIjl�9��z���d����6����z|��d�T�|�����@&��I
#õ���r�q��0OL��H��K@�-��f��NNd՛g��Kl�&��C�ݑ���i3��^<���b�!�m�E�}�(�g
�X#�0�����yL����d�?����];[M� ��i ����S͛�"U	=ʬ� ��	�-��QS����_��M�JQ(e��LѴ��t��$��6���{����؍�V�]�:ᖢ��q5J:��	4����*�![�Y�vl�E�����kYf����p��z���ƈ�2J��3���$��'��W��X%5�ɲkVϫp�*Q�3�6�"c"q�e���9�-~X0�;k�jǣ����[��.�q�Sx	8�m<���;�
�ר��R%Q������G#��.7K;)YX;������uQ�\Gt�A��ݵ���o2թʇ"���ZBۍ/RbW'tD�k�+I�O�	�@�is�3�|ʬ�4�'u"$�E�
O&��Ы"��-�^����N�a�k�#��-�4!
��T��Nx_΀�^�:���6���*�g�e
Sl�?����)�.F�6�O�KJY"��ǡ Iڶ����1�1��2+'��b$q�2���dDw���h�����w�O�z.�7cA{�Џ펫�W� 7�D��
{�oᵭx]uޟ�Mr̂��XMz ��]�~6gB�'.P��[jB
��$�}L���v�}�<e���D�<��R;Ȓ������2*�7�X��de�j�x�底��:
'�$�����D�m��kZ��Lme�-��x����9%��=����I�Q>d�F�(����x��PZW�&�q+o�9��P�f�P^��NH��fiO��w%J��H��V�.�^�N�ڊ	����f��Y`�� &�r�1�Ƀ �RF\���s���~Qq}u���K�8.�_����l��χ�^�C���=��a�{��'�-��A�L2S������!/��#�cB׃==�l`a�3�2~���h+��1�9qE��6}](�<`�&����g�7������xt�5�R���
T ���	E'��~1����& �o��hb��o#�[�1T����Ni¯	�֍,ҥA^0ƅ���l��P�+����v �������~��/���"R�&���3�U�~¯c�$��F�I�3�XQU�뻣��懬�,�9*a�N�W�8������ü���A�Ƈ���	O@鍂	�cަ�zt�{���S�\��On�D�&��!��E���lWG��mQX�a9Kn�����1�j�c��_��$
�"�s�jq��0`�5-��5`�D���Z,Z�2�a�_N�TL�k0)<����>����'�)�-��wK�-��v}z�s��X_�B pb��JAc�+?%�F��~�P`��)���C(��]���4����m)��_2���F4�x�O��Z0=p�Si6�����KM[L�w�e�h����l#��2�0?J�����[z�� ��DyV�CI�θ	$��a!���c��&ջ��P�q�������ƣYB�nv���J���Ȇ�Wcm�_P�M,A#�5�f�k�X)"�W���Ѿ��a�`1߰;�@��w�f��ћ��������jZ-��EB�u�hjhϢt�D�s�r��X�]�o3�O��L3F���u����ݭ`�l7����h#��n�¡;"S��jċjQ���.p�]6�ֳ#_sAvS�u��V{�.��0{�ڀ�"��h�s�}�S��0\x�-�dUi������d�/��L�[d��^��Ye����N�e�.�0���q��y��k�u,n�q1�����p5���ߺ�P��w��AH��؁_���Y��Tw���v4�i�����b�}Z�$r#w��9?��[����l��J侥�3�w��A6�����D����f����F�e���AR�}�w�n���ڱ߁�V�L�%�����ҕ0����c�`���3��C� 8^��{w��]�K��F[�����u�Yl���Ϥ$��<��P��h��&^�O�n���(r�O�)�˦\|j�x��2��!���
:�P��f:�L2��>���	���0�idV
���9m;"1F�ݗ�3fϵE�5��(:C�/�'4�!�$d���N�t��VР�֍XlxVHYEB    fa00    16c0%f%?��}"�b�=H^�F��|4m����,]�lV��NdO�7�據W����Wt8�)��b���Ȼ�(JA�yǤTG%˽;C���y2��ݣ���eK�>H�&*-��i~�7=��e�:�!�5Odʙj��Q��ӓiM2� ���	�����sv�� �sF��aP�fȲ�m���`��G$�I#/8�8�Pˌ�jJ�GX!����[ܦ�n�5�T���R��������0pF��E��HX�I��q��h/TH��~_�oUK׫�Twun,[5��CO��'ڡ�h�ű�0#ߑ�s%��	��x��!H����6i��7��қ`g�o_�)@:G��˺7�V�����<��svf�W��9J-h�W�Zf/ɢ�$�9�v-c�;����P]�q�|�r��OG�Ar�x� ��e��+ԍ�I�Ykq��g(�L�7�cLR��r/ f
wu��­�Ki���?EKf����f���h#0�J����wS�#�r�uw��mt��6��g�l����H��BGV�ܛ�$�+��K��V�Z�����y�ؒ�?���`Ӻg�	]���؁�f��}ߴG���Aތ��$��:b&��ۇ�oF�. '����u������K����s�,�e����d��TC��D_1�������o����0w��[�[��>����LH �ya(�l��>�]3&���sp(�<u��Ie��<��UFA(�M֓�g�+:"��FG-ԽBI����Z���Y�>�O�'/[�Zu�75�$��F�1K��dN�>`�J�k[����͖`��C���ExA�,$��D�0�\��>l�BI^$��9�!����NQ��'Kq׹�#�����4��8�1G�tā�Ɂw��P��К�=oO?	����â��W��uz����Kˎ��f��-���n[Gl���
EUIMS�.�U7�ge�T]�)^˛��#}��_����8N~*��s�������II�A=����n�y�'�k��_�n�f���%/���Tݼ�JQ�s�Kah��Up�!U���	γ��:!�e�ȫi�� �׳[0?h�����#9��l�����6�eg��v��9�=�9s~a�_O�%zR���=���*v����;_,n���-����y秐�t�)�����%X�����Bj��eƋ�(�!�#1�w�Eb.�ٌ����!z�fs��}i�E7y� 6b�-qr }_�`�����M�qK���ϖ~�}2��ڝљ�qI�ᨹt�����A��7����U�;��0��A�Ry>#��b<9q��Ϲ�;1cX(����DK�fI!{��(At�r�kTWa�T�+�O*w�0ȆŒUZ�F�_�����%S"6,������B	�2��x��D�-����sVC/��(ջ.!I0L��!sqv؝�h�)�3��N!�	(
y���ᓓ�/O��Ե۸h�L6�ds�E�Ӎ2�`W��ߕE�G��I��a2�9�}�U6�_��wI���#k�J��3�l�%��WҲgb۶�7��\��^�C�P|
�M_�q[h��q����񥣌��!G��E���_=y��o�s~�S��G�x����r�b��t3=d��?��Lk�P����J�E5E�ұ2�4=��TK�'*ԅF���|�0� �����)�	�&-�9?��0.�c�x�-㐋a���:\���3B���l�="��J嬯*�/���,s��z?�&x�x`������˛赬���3�N�;,��c��ޗ寙�w̲[�r���3)��v=���Y�.r�� �:�*�7w�
�;���C��p%���������t�Z#��M��ϡ���o�$����?j6�ə����E+�6&�["�#o�,q��.��&sJZ2�p~��6h���[*!h/�h����}�B3�̠5���C���f�A�q�@#n�$"��a��G�j�*t����pO�1����|��
}i�fJ�4ykq9,~�wv�;F��b�^��ҚA1����5�Y�d��@��T�h>��f��N�1{Aߴ����[�>`����*`��pNb�.<�"�VE�~@ZT��lp���a�tŁ�G�tqXk���!�ps^���,;�=������tMCW�3�r)*g�,*+x����2���֭m��$+�h�7�jN�>~_y�q<�G�s��wFd�|��!Q�d�+��L;� k4�;`�����@i�%�&W�.��&Q�n�r����]e��f�����vug	)Ďź�|X1�P��-�AE[�d!�ߡ��GrYA6CB�NΗjP���
Z����𘵢^}�xlc�v���B)>%GH�C+1�I�.�}��/��lm�Ut�"yM�#h����둟�ٴ�T�݃/����0<���w�	p�Ѽ�"ͽ/V��5���w�$�W�#��juA&�7+l�O���*5g	�0�����%���JA����s��L�s��v�V�z��&j�7��T����t�����X�QȢ����ז��'u��?+��,��(V��<�D{��E,4*�N�v������:��0-���5(:e]����T�<����J$b8wN
��Ve*$�a+X+s����يAN׌�ל�b� E[�R�$�E�u<��3i���hN�N��N�Ǣ?� |�O����^� ��E󵪡���[�#�Os�-P��N��I�O9��sq��J�f�ۦ����n"�M�%B��^E7ӌPç*1�M�m�{�ݮ�\��邏��٣pJ��3M&���-�-}:�sc��f��J5���T5�3�J�}�-t�!@�-�J�ρm��µ��h���O�ѿ�B�LxkP#��{n[O�ۘm��0"��.�r1�M�gv�l'%���3�|vPc����/��f�s��F�d^o:�}�`�e�rw��^uA��b��x}.X�z�����Չ�N��>�(��$	��W�y]��G��GB"���	��6�4Y�����j �I�[)�́��?�+�O�>���t����d�s�q%T"�H��YL�^���go�/Q)�r��$���	�Ԝnb҃eZ�f��/�i&ā1�傮v�K�$���~��7��SO��G5�*�d��Z�����7 �K"��) �� ��(� �ZHD5F��X�{yk��Y,"�:żձ	�#�V����(�{n��2���$�u)TG���IUʥ	�a�oF�p��vT��\C�8��߮��-bV��OV�H�}k_���:@Rň���V�U�"��z���Ƿ�Ϣ�rE;�&�#p��Slx�(/|���@�Q篪����-��-�M6�ۙ֫��%���ڕ]�i��.C�j3�E�`�:��+vl ��"�k���-��/;�Nl�8N`&"Q����L����Q����5���w�,b�~�F?��/+�	�KOr
�w��6-;�W��L��BWnRS�z�V~�>��~'ju��b����晹p9E���d� " KFI�A⅚S����*���_+.�ƹŧ���1� �)�(����u�biݣn8z�~���B�S���8��0�UG.���϶�4��vWE�����WZ:	�snltB
�j$cy���کhh){M���(@J�fZ�2_}wn�~o+��>�;�j|��0\��������e�}6�5?��8[�}ށ�̻���	B{�,\h.��\D��BE$��92�;����y�1�?��,7ߛX��)	q*��Ù����ZC�v�?ٔݦ��j�S��h���������]��'I�?�wrc��$��U�K&�3��V^}���
��(�N�e=�i��-��G�4͆�Z!M�jZ� �6��_2����>!��"�2o�N������PҦq���K&E���oCH�"h�Yi�s@*M���,\�_`�t8�9��eƖ@�K�H����w�ᘭ�1�k���>�����h�5S��/q�m����В%´���B��I�Y����s�e��&������Z0�����PD��m��L&!�"����kp��+�ڲ���k�d��W���$D�'�\ֲ������m����;DH�J��Ð��p��5�9=%O4���^�����?�)``�/��u� yL�R7?�vq�lѲ�X�"���L�CHB~�m�5nZe�M��$j{��NY�\�b�	SY ~����A�n#T�ӷ�-|mk���'�/��^�6�Tl9�D�U�1ܪ��NM�MB2����\!D��i*�Q���.M���٥�L��?�ECf�&:W��' ��y�S�++�U����:3�5����/gz�㖊N��b9�\�*�is�7�b��pܽ�꟠������-Xb�Hׄ��=���rd������eid�Ʌgz�C�d�|#��QX���_����>�k�b�[�\�wͰb�PU�И+;��Ht5b�Yp�K�K���M�`�l�LTI�|n�F�]�!G]����e^��;}�0
e$����N��e�Z�=�ݵ�}G���������<&d[Eˢr���$h�l�0���*�r~�C.�npko��Wf�f�����Y]��(��@hil��8
غHN��.)7=� �=L��u����a/�ǽHX��=�yy�p���mp�vxʛ��j�S;��V�$\���_��r$��='���!��X9��85�_)!+�G��`gN+�;�B(��;�D��Z&ާ�u�h��b��N^���eP�#�	����(M0S��[���cԣ��GG�/�*��hf� ZhbP�E�3�%���a�%�ϝ?����-I̺���r�qe�}��X��Ol]��������$j�=��h!�?|�� ��#[7+��a��jӶs�g��x���V[��w#p�sn��Y��Ā�p���˕ԍ�	B0ļ��@6����|�3�^��ȚG^t���܋xa!����0�4�F ]J���vԖ��ᣀa..��e�T�w�pg�{���_T����>%�L�b���a˒����.łOƪ���ԲH���̑�?����m	���5St��i��`~��q2#���c�Ǽ��<x5]L��TU�x�gD�I�qA����n8�{}�e�5�z�)?!�<�����v�6.����f>U�"$�j�Z�E��R��� T�&LUx�Eq�����؀���.�ՈG����Q^���8F��-���ǳ������R�B�W�w����5x)촊-E��y(�;��ʵZ/���A����>���kV2�4l�炶v�n�[�Enf�W?�Z#��:S��z��؛$���A��v*��8<{#<�
o@���� m@��/"�i�y��uSFVZ��IL]�9�FT�d��_�P��.d~O�Nk������D�C<K�=� %����kb����w�B����q+B
]���0�p�]��o��ɟ������9V~R���
Pey�	|u�:"�LP�n����_�̋T(OD	�:��N�)�L�ibxx����Br��V�`9d��r���zjW�D��F�l�Gw�$.Ub}״̇����A'�hH'cߵ��"��2a��hM@��'7d��N��%�v��G����88i*�%��U�K�nu��1���jy�����W��m��������J)���S��H�6�A��KQ�cԭ�����u.�޸�,���r��q���NH��:F�w�z3q�V_��h�=���-�TXlxVHYEB    fa00    1740�(�J�Ti��>$���nQ���x�lM��4X�,��Z�3u*�47>��BCzB�]����ZYbn�jH!~W
�\�nL�*��Gf
������uU�,m��W�j6~��k�C]k�@�xy4����a%�I�$d��d^�"��2�c�W���� ���'��у���L�_����kvm��Ԃ��Ś�-��4��t��`�?~��D:�9�2�uf)�JX�w<	�\
�$��7:�k䞻Ѫ�B��zWj��HV��Q�L7���eU�U-�n�8�w,��	)���x��FV~;�f
vO%B��cZJ		ٚp��Ǘ�ӵIU��B?5��8q���7̂�_\�f�!�E���¡��9їk�| ư+!��<�4)��j�l7���z�G�oT3�әu��db�3��ɾ���S�foZ���kxQ�[�yTk����c}�u�iH	�<+s��yH�w;=�,���吲(���2~���݅���,��b)���5�¢�_����Kw�h[����&4��_U@~3G����,������8F��O�M]�ߣ0F������F>�`��DN~��o�/��*c=��v����'�������ݮ�E�>?��̚Z�^�ʘ_~�ռ�Td,V{��g8�8�i5''�wq��!&$��c�z�	��Bw����m���b��N<N�
���!���@7�PP�`d���>�2��"��v�4��O���x��1w����>i�ې%��o�捎ކ}��9{�p�6@��%ڊZV�qP�Vޤwp~S�+��VT�y-9ж���M��ބ5��5��,:-)�e��?Vi� �}���S%+vp�g5Rf��4��X+�Y�F"��z0���J�^!x��s�==z�/�/�J�^GeDEb`�샟(P���(�!�8�jVZ:��^޷:f�ZR�j�- ����bM�3�Avs�z*���S�T}.�$���-n�Ӷ��j;8��/��I�$�|�m7t|U��`������*�Y�����:1�д��1�<ݝ�,����^�n��P㞎�&�%)8��r��k��22�٣5�5$u��iyE��@��VJ�k���9�,���F�MCU$��f��ÑZ|��.��}��lU�JJ�/�])8{�Xpy���L�qw�Η�jE7l�Q�tE1Tb0k���e�uH�Y���9's�i)�ۀ��S� ǢuLX�ʎY�dG�_3�,����)����ߟ�ӝp�y�g?m��>�uN��p��!����֍�0/�a�GǞ�/1���~�Cu�[N��E�Wg믓���h yQ!	?�KL���L:�e�_�)i�V��O���uH��D����ˣ"�^���LA�M�S�p-��:V��.ta��t
�,J8)��\([�	��ʥ#�oTmԣK��2K�^-~�j�.��*+�Lpi�~������J��ƗD�C��
�M���E��,��%�͘�1eQ�����XX�B�>�.�e	r�3|$�Jn�v�J�A��T����K���B4��@�A�����o���w*��-�Ӌ���?�.�{�;�[f$r���Af����+�փ�gE �$�1��A'N>A
��o��Kv���z����(�g��fU���,���;�'B���ax����6������[M7	1}=�	fK�eH�AU�1�� �Ӗ���,-�bՉ�2w��KlQ��[P��G�[����R�>T�5���0O����E��"4�S��9~:{{~a��5�����$��rce��\�1�ٿ0�Ď����(���u�>�l�
#�Ӥ��v<�0Ӗ1����*X�AO��Q;��4X꧱_�1̵�r@P�*È�to=ce����{������JM�=,jF�����hI�`w*�z�{��ǐ�w+�y�.��3v��]�Jv�-�3a,�e�q�E�Nq��?� ��&?�P�s;�����+?������x�'���Zj����v�҉O_��#�_ei��l���Hf�:E��H60��tV���	י)_sn�����z��.�m�3���^4ݴn��67��OG�12"B'iێ���˵����`C�Є�F��k��>M|n)���g��.箕i�'/	d����tbM�k�t7k�Љ�1c#Z!J���|�<����^�c#TαXS�(�1`�E$�Q��2��h#�y��:�M'��牨.��|V
��GgF5d9j��g�ʭ���%;вP:��3H>Hcq��"��1������`w��щ9/ZY�=	�&��Y%3�Ї"�ޡ$
�������`�z��w��O���Rף_�r qeJ�$Fb}��Z�~]l�F��o����kN�n��NBMW���=E�Ĕ��z����)�}�P�ĝ<
��������t�b�GGL�C�������R�(�݉m�0�
���A�̱��[�1R1�p�m����bx���E�8��.1l��~��?ަV~R����d
�����í�ĕ�ԣ��~5y���X��@��b�dy�D�5���S_�՛b��t�Uu�S����{��A���j�ؘ����V:D���N"�H7��W���Q��zx��f�G��%��̜����%����}��jK���|��N�r�����!ɀ���%��]����6����E)C��4j���y��Z:�ؔR��|����V4W�SFcO�.�Jd\&+���P-��_��p�����B�E��l��Dj�r_�C�j�Mx%RІ{�7강A��Bz��O����؊�_�'��׺Uq�Z�{��<T��~ǻ'B�u V�(��J�oZ$�s�c\>��d�/���N�@k���HTfv��}�+��ƙ���D���c�ؑ�ù��*�2ȇ�%�C����C�Z��ke���`��2���v]����]kOU����J%]���6_#@�M��՟JR��c�!6!����x���q�]C��@i�E�o�|A�	�Q �k}���w�D-�"�*/�XNP�)���x������Ψ���+*�v�'X���q��թ��rմ�k��(��ަ�
~7�X�_�mJ8zO=YG9^L;0텥����$3.�L~t:��˕	�'�#.���->7}�G(QR%r�$�7�?Z$!3�ڼ�ז���h
����`�cc�ܫ����^\���׼��}�X@/T��̬��)yZ�Һ�lm�#�4A?���-2OF/�%�-�c����'C�(����B���?8�i'Ӟg�W���Cgn-9�{���u�k��[I������U�����ՌMp�|��
�l:٧kbc��q�Y��� o߭QѪ�el��c��QI�.�ω+�mA*D�۶�G���$���4`�e4S-&���U��V�4�)U�+�m5��$��PՂ��W��ȳ��H�;�~;��Z{�B
�I1��%:�hl������,�?�زG�~<�D-�x[#�t���G��2�k˂
�CH�c�A���Ǿ���S�W![�G�����Ca(�G�O˧Aj+{��b4�m�����A�*�[�@�R*��Ǣ)�c>@��&J��!a��N�����b4F���wZ����v�44�ִu�8-�.l3/�ۥ�b�H߹"%TZ�9�����	&�P�O�2̕���/�`X��c��\�4�f�}���b� Mn-$Ae̩�>��RW4�7�x�
����쾀#x����5j@�i��\ù�
�Åx㝸��̺���c��9�
yaIl8#2�|��O������8f؁5�����(<�D=nN�nݡa������f��e��p�	�{�Z�c�����������h2T0����$�`��52<����zc��W�,��3����_,�H�e�Y�I>�(�g��}��W�j�U'�mMجyה ]6~I�4:�#�>�ĳ���b}g/�5�r�ޕ���d����/q��){9�
�:[�!�9�j)x0*�G��k��t�x�{�%O�&�f��o?�B�`M鬷�ʿ����(�U7}�:d�j~cv�о�PN��Q��r�b���
so�#�P_{��cԐ��݄pğ��]�×���j�4��Y�gXڦjj5�v�܈���!F�����zL�y�W�Aa������,G�i#�-��E�8�/A(!I��@a��:�Oɵ��ݿ��8�Xm6QLZ4ɔX���z��C�M��t�Rn�Mb��>��ZQ�3�I�G��V�`v�u��>G8;��'���nwXAf
KGw.�Fd�� �#0��:׆w������t���P��MI�V���gU����u����lq0e!�"O)�;��4���GC�B�(���Y!&��{-ͅ:�j�M��DK`�lՙ_/�
ڒ�19��^���c�j���~>�Ѻa�f+^$��T� q��)��á�u���9E��-�-���zJ�4!�\���Z��,T���i���*"v�x�]G!�@���ZU;Fv�Ď�g�Կf~6�y�Bl0�H��8A�U�����e��S�
�w������ou��a�����)��y���Lխ�F���f3�}V�aQ:a_"��15�0��M�h��lw�6�m}s(���r %F#�J�I���y�,�ʓ�n��U�0~�	�i��&țhɃ����6V�2H��p�ث�����Z��̫�ބ��8X`������(�ǧ!5>"|gP���N�֋���pmo����9���R������I���4�@���$�,�+,��n%��/�U4'~��97����&�����VKU�	Y���k�	�B�˷��,��c@�y1t+O�ƍ�>�r���^]�`Zfv��eH4q�BD�l�#e����й���%˺_������{:*�&�*��m�W@�dvh\���?�XV�8��E���ו[鴒kG��Ø����������+�a�I�Q�G�q���{{W����I��^ZI�����
��C�~�<��<���1&B#�������ړ �~f/��ňr�}3^�<s���Xm�p `��	��2��z���O{.�}nZU��@� �.6��d=�tJ�e��j��|���n1��"Si0��/}Gw1O:��C��Ú_��;��a�h:;��M0�\��<w^G���a�Z��j�C�o������Ց�m]��$�4H����r�x�7J�=��aFw�y>����]�^�?�|����L��T'�|�)������`Ҟ�@��P�M��6ķ*�������<r^t�S7��d��6/� ����c�z<P���� ���ymh�Nۅ�#ʎ��M��q�p��I��������W�JK��� <�h~���������p�AZ�W���좈��2�����[����Dp�E"3f�~��6���n�nazsi���VRA��v?�&��B����g?���� �Y�:��ѳB
�Sb�����6�G�����:R�#��/�kRj�$�p��`'����}l����+mI��@/&�gX�U/�?�g�r4��?�x!.?rX�)�2:H�"��������hG>m�}��������������O���@�@�[�%��c��/��X�"�PV�����O���eE*ڄ�PiqD��m�i��$խL�D�9�uz�Ф,k��6�o���.���Hl�"�ҡ &�H"�SF���|jV���ҳ�B�Z�(���x�	�G2��Z-5�P���
�d(c����-u�Q����&N�q�z���N��������ӣ�>n�%���|�Y|G.<��w?��k�����$�NyBi��e�R�B�ID�ͻ�߾�=�
@�aߒ��*_���Tx�}�����1�	���-�m�^���XlxVHYEB    bf14     c60�L)g	�x���{�i����>g#I^�|J0ź<�`�M�P+�;� a��nX���=�t����<M�b	�J凴���B�Tx�������s�T��G�f ��+ڟ��7��(��w;U��Ɛ�~�l�(�У���'LJ�Q�b�?>�#�� ��%J����E�oy5*����&"�����z��^#2ڄ���oli����DT�
Z�T��2�kQ6N�Y�����R4���FO�u.����a#\�
�ڙV�mnk��$�c�E�(���č)��
��F��V]Ci�Kv+��9pA$�&@z�H�S,�+����6�"�U���a��x�$	�V��Y[=^@�B��4w�dYZ5�E|���`��lh�9��KP���lP�)w!��d�6��4�MN���󧧠���ҜUxLP�3^2�_I�İQ�����s2��C���d&6PQJ8�X�˒K�~����9��r	N!`�8X/%Oy�,U���"��lb�C&����8�x��M
gL�鵬q����ۺTMx����OS����&J�O3E����S��#�������=�����٩�& �ǵ����(��"�D�e�/������gp*Ϸ�K�٧:����ڱd5�MJ�-���	�u���U���il�.g���rv��0>��:�Ϻim$y�_��Vy4#�����c(���)�;��&X�d��ٕ  !FBzI��LkY�Y����H0��h� ��&�z;a�{j̑��*[f��KH4��1�s��
wհxh����+R����OL�At�5|S�.F:�����-}�?����~�}��O��
�O�����[��@{���p���U��4��pz�0B����L���CA�?���f��v �҃.ܥ�b^)kOTI�M�V��A׌C��ڑ@�j�����7�h�Q�6Q��I�n�Q�iS����"����dx�����J�IH�O�7��3����l�W	C,G%\���Tˇ�D��,����ȾL{�i2])�^��>2�k�!�lo��G�>
p�Q���f:1��M�"���+�b)��SvQ�q�4�����~��]k�M�\Ǧ��}L�t�F����P{i��O��l�v����K�Q��8�MB�qe��W��b�K.4G�^�۲K��k��	x����X�P;5�< /�,��uAF��d
զ�q���.z�@��e+����9��su#�W	TG�I�wyI�\�_�Z0�3�.�3�Dd��,[z�i�`�.]�w���e��v��$-=_��WS��	�����~�ٛ�J�tiv&���"�xo����l�"Mړ���dx7!Q��<I��w@HEu�3ƥ]�/<˾���edl��-��=�7t�iS6|�"J4�IpJ�\^�-i���*"Wc�����ܸ�8�l/_��Q���?���S��ĭu���i��oh��K'���:�]9�5�ޟ���b�!��^S馪t��0�˅i���T���X��5N����d�̭�1_
i*��T�>���}�M@���$�F�� y��%���W�1���~��:JA��)u'uY��q�º�����j7�̔��7����H�h*2.9A,��u�/� P��=cÏ��*=����1�x=�2"0Y=�Y�J���0���2p��&�]<^����p��Q��ģ�WG;�8�v5�e�U��iFU�c&y����6�h��V���<�{����x#��c����[2f��ha��/Cl��O����A�;�T�,�đ��!���ݕ:�1���F�}Y�FQ�VJj�O���]^��3% d&���Vv�Q� �G,���4����4�=nv)g^�N� �5�/��F�����%4�nA�Y�O:�����Rr����4j�9��,��#�+�"<G�Q��ق;�:�E��6P�������Y��D�,����1�Or#�O$�N�)8�ALi��'�s��O�7p�2��o�ɆA�0�ĸ�<���LV�rv8l�0��S�*WI�Ұ��n��S��X�F�G�nb�Q��luz\
B����.�9�{���K��T�IU�����2�V{J��bS	�������(aZM�	ކ��T\�lq�ܷ�cR$��'|�gb2K�{k	�sa�i]�D����,{������Y�[b�*�ϭ���O��5��rH�M�pL'i��
��/�C�����4�[ �z�_ 8��#�8I3Ht�:h��~r���*�C��``|�n~�X��jE�/&&��֓�h�ق� ϑt�<.ߧ6� T��9�f2ZJ�2U�n�jn�' ;��J)T��[�ї���o�~�,�h�m�6h�j^���f�-<�E=�c��tp�W$|=>�?������������F5��"t�;~�����se	{��F_XT�u+^���}��6�ἐ_Ӿa�^�+������R�A�m�K�}�E3ˈ��~ �a���ܫ�ץ��2��vvF)F&���(K\�7�4m[�RSd
�
�n���=F��/biz�L��!L��"348Z�i����P���g�c#� d��L��zt���w�eg!kV���80IV�kI��"�|�|�j8���v������J=��Xx����C����!�{]�|�	��wa;ӂn�+�	T�Ӟ\��5LV`�E�_���_+��Z��:�4�?� 4��K�~aY!�wj�B�k�rq�q�y���y�OΤ��ꦪ(��d���S.?�(Ɋ��uV��H'br��f�T�>���f(-���oL�����fy��L�j��I��2�a��&�,8IU��3wk�jl��A�B&�QK���ݺo����"o)��|�z������\j�j��0�K}�&�u��ѭ�@n�?��B����v�i����|#>�q�p.�Gٴ^̸�p��{���L/��ͬ�X}���Ϲ���KXd5ߣ���y�I�q����42���E��2o��L_�Y����H*50�=0V pU�U8�CKH���C�4�Doޭ���g�O�,�-?}a8ܗ�`��H��?[<U���YZ�ƀ"l1��#����+l�4��4�L\�>�})ng����[d�$���S�07�X?;t�