XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ރO���2wA���oH���]�TD[̞D�e��z�2&h
���9ʂ�<���$���DG��>`�~�'.��+M��^�`ʨ^�1�UVD�j�HI���I��%�.�F)�i��!��(��p���%��B+��?��8[%�ylgDĘx���h���({$���&�B��ڂ~���_$��g���\2�������2��E�5=��ϗ�۪���蟟�ߤ����ژP�A [1ˌ�c&U4��`�[v��.^�h�#�*��3!�U��5�j)@���ï�r$�t�9��5�	\���H�����0��gN@[�fI��������� [!�!�ò5z�"OF��R0�g�&6��+�^�Q/+@o�i�?�O���OR�hi���fC����R�B�&!p,�u���.�mu�~z�O�F�����:��w��J���y�Ek���h��	�ʤ�}���V�^t���0J)��m��A��&�f3��(�����qx����[;�� �B�y;e�r#q����F}�!�c�7�2K��h� ~ˤ\�j�U}��-�i	>A��^��51��p�H�[f����'ڌwI��^�DA�UФ;���ā�,�V��2jB���0���&��BW���
��#`�9Om< ��Tjd�+�]'�覬����*�����n֗��|���S�1��ђ��M:�y�#C�қ�Ox�X�%��J0��)�,���l���%��;��֓��Ɯ��Y�Y��^je����^��XlxVHYEB    b8a6    1ac0�:�l}q0EK���Z�b�<�؉�;OdG(��>g��qľ�9�>.K/"��# �6Z~02:��g5�mbM(��z+�:$S='������%��UtWxG�h��\1Q�]jC�J��۩/������Ezu
kÂ2ax~����Y��ő2�h��)1����`
���@����ȥX���~9@�n��4��R]������2K~��9�����8_�5 &a�Q�C���MS$4��L��ۤ�d��6S�h?���H������ZW�Zzw�J톿�wڅģfc߮��n��β�-c�⟺��N�9�<f�Y2�<�W�CU�Y|�E�ES�ku�PcR[A 5z��4ᔚ���}��2Q�8+Y$]�*�tvF"�\߫ن��(l6fH�6�M*���k��*hnfq05z0��t�d/L�M�I	M��~�����Y�#A<�_�y5(9B
��[OEّTV)m!�
�+a�`Rh���S���@ Y� z[/�ˏ�Ϥ扸;u8��E���~��S�t=�9s���t�1RS%�2�*�غg�$����>�$H��	�D�4��T��Bb�o?�����T$����.��>ͺ&��}0���2q>�����v�+��[�n��� t��-?0���3�(�=["Y������R����%̪��CD�ċ/ϯ2sk�_��<R[$n�[��l�A>�p��u����#��_*$M��l�iiQdx8��b��ٙն�@o,�-֬Y�M���A#<_:��F/��M��\�S����h�%j|j6�9� �vsw�@�׀��0���G{�IIS1�W�A��sx���B�`{ 1�2}���5R��1���ZLUk����!���B;��U�v�\=����Qvr].e���:���L�B�CM��Om��0:���BiJ9�_�;�������a�vu��Wg�����z�~��Ī�3p��h�|
�g<�P����A��֙K���Y';�J	�F����w���� �v�x���?n`hz�?���{>IP�*���^-࿍ �\�b�K�*X"��2P$8�߳� Bd��x\A,�F&8�U��L����_f�z|��A����9:}֩��k yF�2��svTSѧ΄�Nכ�s�W�6i:�L�|,ߣ��ݨ�(�zmr�\ôl<B�u)@��d����p��r�s)�7��S��2��U˚����}��V�y{S*џ�"x�Q����Jc޻��0=8N]d�7��]H�j��k�{���L;F!I бyJ�@a����bi�)L
�t�^�qݚ0[�E��7��x2Ǜ;�&��q\I�p���E` ����6i�l���*��b�W���l"G�ֽE����M���8��
�+�~8DM�`�~�O4`(:��A;4����V��\�\X��@����Au�x}I������7%Z�8%O#�2��P�7����^ ���)�%�R��)��B�[��Z�*5q?�:�u[�9�����LzW�2��&9X쉚�;&RQ >_ܱ��D�2?�`V���}s_L>R���4F�r���3�z�)z4 �I"�hѶ�刯�
!&Kh:�����{j-��n�J�PğW�''{�A[�1HES����F͊�h錹�.@T������a���	�q��B#�||N��Ŀ�h4�jD�%2׽�R��U�bOQ�6�c����ٟ�r��Ǌ��{d��?���� �d���̢pC�S�Y�D�j�Ma��(�o�'�Iu>�fv�qj����*�+4�%H��Cb?������[��F���.��X��Kw���eМ����Ik��J�Ƶ����9�����Z�+ڒ+��y����o�F��,Ź.}�c;��;a0p9�J�[��UZ�Z�t̋����H��^��<�la���0B,��:��rU3�~~%G����R���i���!b
�����
e\�W��u�5YN������W�
�~!��o)(G� �Ckw�e�
id4F�ۑ�t�-��j�H��&[M�V�s�,ő�J���726��i;ł-���8:a~RPT�\�<Vi������N�%Gx[I�֛��zv��v��N&:��?����7�"C���LR�fE5A_�k�X���Y����*��l�Yu���$ZCn�,�b����i0n��szV��������8�X�a��P�Y�l�q;rq�!(��� �r`�|��cM�����]6A:G ָ`<Ku�fb�Jm#Y0�!gI�v\���ozXaA���1�z��<�D�>|ڕ\40�ݖa�ڛOm%�&		7��&*��~O��5Xҹ�n^ʖc �9��cyM���=��u���:~���:~.��|��ǜ�H���M���|�{��mY����\��*���6B`8�R�K;����n��]ϻ�G�c^�Vą�\���ZN�.Σ�X��d?Z�M�J��W�Q1��1;�ˤ(�h��O��'b?���XBz׋;�b"�%��a�q`��S�bs-e�������0���G�b'�~z�$慇�*kG����l�I�<ʮ7����L��ν�g�ߑ��A�ڪb�|��D`� ���cm_�UyK_�'�`�x���������z��9�j���TL��ND���p� �o^��X���My����I�7���u����`�6[b�x�>�(#��P`kD����C�m'[� ��ijW��x٣�����l�+��}+�1�V�n,a�P�$1��Y����L�_�u#�3ˍ���R8��s�������z���.o���&<3����Q̗�:F�n�ҋG0�!���s���C38�h�a���$�N�6Y=VU�^'��:�d�2�5��z�d�f��5��0-�]���Q�L�����%�Yv�2�|E��3:�yV�S���-�����m9x!�gD"��R��\�� �����Dv|���&PӺV�Ss	�y&��&;��͵lV�[(��c������m}�2�3O�9$�* 	""�ڰ��8�1��%��S�/��sP��}wP ���{ߓ�-&J��xR~���jd*���z`���a����j��T.�Z�Г%Q&���H�T=S�љD�9���t�z��2�{��D���{>�֐��BPؗ"�B�d���]������<���u�J��]��V�g�z���.�K?��Tg�z��[e�2�2���l��	~vYo��Nm� ��Gu��~��\�� !�����Nw��AW�e��K�~ҷ6����<��I~�$�����U���1�ƅ{��s��V�tp��Zzr��)\!�Ɠ��k?�7����f�k���`���ƺr�:I�9:�Ts�ۆ��<�c2cBU����|��ƺ�#U&�C��mt�G����B�헴�r���`z�,z�/6���	����D�oM�Q��d�d�|��i#�z��c^��[����v��&����~���9��v�'P��\O�[]t����w�����bM0Jv0С��H�
�:"�V�3���	�\b%8�^���]X=�~�C�J�A�IN��jk��H@�M�&���ףu1�dA�ŬNTãܮi�����3����`�'�V.���3'�f��f���g+��V�^a�n�(ȩ�'����5�
m��Ds�#���@0H�O�oW��4��۔K g/ُ���.b�Vu0MD���g��=-*��b�e�N���0�6���k�ώ��v�mm{�bt��p�ڹg �/P��Is��+N!��m�WT�r�ߣCQL��qXZ��.F�I������4���݂#�� ���)<�����δN�ώ�fC:^�O�s�=�Bv���Zr��~�V�~�΀x�{�XR�<}EU�YY�i-�����&R����S�|P�J� o)�t�H�O���&�VI݀�$hBY�NP0�I��R�`�
`�j6��w��������x�b�/�[%�NnKЭ$t�0�˽ 	=�3ЦJ/8d�Ǳ�1Lļ#�ƶ��&پ�ۨ빥_��l� �ݞ���Vy<FR�b�����M6���2zOW�~���8c��h�!G�%�~���D'鈭B��k�)�;0�6��b��Y�4Ŧ���r�D�2|:�9y�|ч)=Edf��m��3�ڙiqDt-�l�����5�'�����gU���ʀ��p�t��C���q6���<ƅ:n���д	;g&��O8{�e��������,�C]��'8��'������4 �?kn��0���l5 f2óάw O殯Y���'O���鋰K�߶+�Q�i�n�{���-
�ҋ��v���a��z���cl��d�H�g���Ŋ����CBȓ���@���ԉ�q�꛰Iy�6qǭ21��U���d�ѥf��)���F�� (��Ƿ�AD�џ��:F��-ڒ����n�$�.`.��WC2���N���}*nc}�J1��v>�fs��,/j{�mسO����KcAR0�3}��,��B:-,�l��D{�W]9�Wn�3�cϭ�VbH�P�>���Ǉ�6?�ԛ=�[��P����D����k=�sp �I_"��PZvzr "���]�2��z)��C�ǻ���_���w�J��rT%Le��]��kt������25IU͢��"$I���j�!F��I#����*�������x�Q���ʕ�[���h��dd�0�ڽ` !P=�if>��kѕ
�PU�m��Bj8��1ɕW���]]���4xŶ�W)����sPYp@�g�1�;lK���9��!u"�e��wP.�y�{��Ը�f�x �y�aq@�vU�s��3����P���كrn�݁�Ùi>�����\^�ڗ�vۘwl��@��["�bwc/�.�=�6�����ٕ�Ҷ�:w�^�o����Z����X�$����m&8��K毲���\�x�lqb{���y�|Žg�2M���́	g�s[�r������T�U���p�WUӝ̮�k<B�F^�1+P\L�s4cL��c+����Bo@<��B�Q�0;t��/����wlPiF��dص� S4\����z��n�^����D_��vuKY�oޗ���K�y�ý.�$zY�T��n�V�t��W�)k艴�	��N�݃+��6k|v��*���OH����=�q�
�)T�v��($_y׺Fs�}��tU�v/?�o������G�$����TF�w�/W�Q�(m�&Ā���T�1����NZ�i��Q��7�nR�[Gц�k_�l�^��s�s�_Hv^�_\���U<�H�@K<RǷ��*X����4ea�k���W���A[�����s}����%�(��vI/߳�[?J=ZVZ��2ڢ	=����jc"�8c��o'�����&� b��g��{v-շ�q�5{U ZŎn���kGb�_�Z�6D9?+:���瘝����v������� t�K(�;�D�_�Q�8٤.M-!��tz2� �P]]�7It�(~��{��e(	1 ��~2�׋ͼk6(�*�3X�Z�5q�ڙf��+Ac��|2���ˀ*�t��J��E$�(�x)Z�gY��S����W��� ����4�|=-awES�\�҆ISN��QM~�G��˻[��W>�3�:���~���}�k�dN4����m��ގ���4,o�?��~Jm3�VKr8��a����Pl Mג?��D����k��L�~m*e�#����E�� ���wi�l���K��Ù�j�^m|�  &��:�!b^h�)�ج*Z��\�?�G�┆C*G	�ĉX=���:Q�����E�4��$t�̢�1�Ɇ��޾W�T�Wp�A$o�6�W�e��m��@�Y��a2���v rK��q�[5�T�MkG��"�eJ�3w_���HZpIo*�w*}�eV�KU\���������A��o��
z��x�i`de�eU�$]A��2�<�G��xx���D]�c�WX4�݃6�-(̝�ejE��3�>6��K�C��h��ص��;�/�R�^P0qq4��7�����g��� ����ʝ�B�։J*�����O�9k�>��������)��6�����|�Q�����x�v^f:4GC�.V�_T�sy�C� ���b=�.' ԓ��-Gl�*���M��$�&=T�<��~T��W����6:����]P�_��W���F�� "Z��֡#�e8���.ͦ����u�(��Q�����\�ߙ�Dy*�\_�D(���gMV+�i��m=�w��cU n�f4���;��E�|�u\�H�PTCp)9�|݆$�%d����x�`rLju�f�a���r8c�c��|-��7A�Xlu0&���:�Ε���P�1��%b�6R�PjRZ�#���X���]��h�:_N1�FӊT!�������V�^ʥ���Ƌ��1Nf�ض{Y }��A��Sb�e`BS�Θ��ڐ&���:��0��w}�����Bb�S_��<-:MI[��|P�+��2\��^����\�S?k�|�rU��2[y��?%8���O���=r�+?�N�p\� ״�` E��r��fc���ܶ�:A���Q��8'M�4�F��-��T���2�z�d��Mx�����}2f�,V?���l�s��>��W�}ų7#W+J%b2V�u��ˡ�s�