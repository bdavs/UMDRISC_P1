XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�o>y��Z�]��������Ϩt*fpXqL�uup(�*ȉg�"��Oo��
`�&0���>G}�$_Ż�{�A'N�-$��s&�O�6j�Ǎ5U�dcX�Q���H�]
�=����ͧ��b1��U\8�L'-��K]�\�\��P�^i�v������Yᘬ]J���Uo�j7�G�l�3p� �V��%��[ez'\�Ca�����:Z_}�n7w�+BĲ����o�@�o�k{��C����}���\E�	h?%��Y��m��,�P�B���g�%�%�Q�YQ�l)���|�����4���d���(F/�b�f�k���BR~ƪ�@)�SM��K^�/E�A�E� *m�gy��㚵�_���;��h�g���7�NO.����Q�y�>L���a?G�z�`l�랷���Y��1�}�Հ���f+Phf�����c�Q����g��UMؐ՜�wҜ�=hZH��y7�x�����{�g�-��,2���K�a~ |���ӷ9�A�.d~���o�\��5j�^�x0]�Oד�7ex��}��������v�a��Q�J��4H���|aYE� ��R_d@q5��/�B}(�������R����6��|N梔I;����s�(LN�� ����>Ay�X�6DC~ԍ6 ��	۴[h����9��Qm,`#Ե�Eh^l��@os����$Td�̜c2�ܙ*)��n���Wy�5���[y7D]���0DωQ1�XlxVHYEB    162c     850�p�g	��%�=��ϊ�>����B��K���}3i����h6�.c��i/�q�|��H#��;�W����)�H��2�w��d����:_��CU2�A�_PN&<�Y�7��͡ѳ�Dl��Q@���둮* &��	�°}Z�3�9@�����fߥP�����q_��k)n\^!nt��kOU��9򰃚�aFZ���n2�l߱�il���?6��aҳ\Ws�}	5C��Ï(-�ܦ�Կ�Q�����JR�6>�,���M���3 ��<�V/8]��o�C�+�l4
���F�ꨇ2;x���+�H`N=�U7�w�uZ*���]@]"#����37YA� �,Tǟ"��y/��$7J�bbG�G����G�q��D�Z�2�AJ�^���|w_�[S����+{^|U��z)�{ Ӫ�3DX���jhbi3�6u8�
%�P=��t��c���^rw!#
�q����? ��f������+�w�p�&W��}�ɂ��6���M�j����b|J���;���0)�l��Iݠ�#�UH�ؑ�(�v1�8x�pz�1�P���U�I�%nS�<o��S��N��H7����-�DT�Mc��d��i<Ì%�vk�Xm��.��"�,�����ߥ��?ߋ��Z(�o�7f���ܼ=M��WMo1��'b5��R����35��s�+���@��p��Y��}w�'ҍ���=V�F��Ф�wj��H�	=�l�P��ڎ�%�xp	T�������d�(�q$��=��[���\��~5Z�t�s�M��D��9�V=/���{�M�i\�_>�߬�#�U��h���8_�"<Qr�+v����v*��T9JbJ���$�E�ذ�!1��/fm��Qc�݉�H�9��*���8RQ�e|��U��д�?�'��ͼ�z�Z}H�$zb�
C|�K]|z�[��3?�g~=�~pL�������8
:+	�U#�ٺ+�
�V��
L-Q���N]5���M�P���6��H���������^��~(�G,_�
n��>�lv��V�Q�i��w3�T��/�1*\@�#�(ۍ[al��Ot���iR�#U�����k�~f�%s!�|rj�-��0���>L����J;�|������I�}�W=���ᡀ@��y� �)8I�yÃ����*�},��)��o���ďs�\�=^N��g���g�N��/'B�i��{?-W���y;���ˡ�f���Z4�\Rӄ,��B�Hr�7�	 �!{��Z�����C�V��gQ! %� �X��P9���$-/�?JM�q��_���^k+�ʦ#c�<BJ�k^*��F�u����oԺ�rj��3O�e��Uy>�S*5 {M,`ͧ�v��`=������N'�����q��e��2�����A_���_լ��ճ�������a*\�.a5��F��AE$f wʝ��/�A�7�Qk��¡���z��h�gZ��9"8͌�0�	vW���ڒ;K4��GC/�����hl�����<�V�7��=�*��ʔ	��	�<9���TL�ԈS�#Ϩ]���j�~��gq��r��������ɨ�è��&���TD��0�ȱu�^��\��8�/�}k���^�ѫ�;wZTzz-@�2y GmJ�#l���'���f�IBDX.d�'2h��[�Un�&*2��L�Q�w�٬a�p�xFv'�����Zs���|�m@R�Z� &�*>���-��4��xtC#��Xn X�;�8���0]�����g#Փ�IA,Y"鬔^�Ӝ���H�{�s�R�"՞��W�@�UpP��ʓ�F����'7�������:���zR/�Aj�Ӫ�K)>�����j��Wg� ��g�FGӐ�5���ӕ<���Dx�AO5٣2��m�� ;�	
����#	R�V�R�$<j�çKui��6��D�Þ5cI>j��r�(~_���24	&��?���?������U1B�?Cڅ����E�B3_.������p�ACo��>#o�-{��j���i�P���þ�Q�64P�UD�o��{t��d�"M�Jɵz�'J�����՘A�I�����