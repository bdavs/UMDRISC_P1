XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����N�m�x�Tם\�a�D?�߇\3����`b�:�+��i2'���&�ҳ#|'�5F=�C�iƔ�;��խ��X�'���fW�Ā%L�na�d^[7�#GoBq��{	=@��PzIVQk/�EuZ�|�����8j��2��a��˥����I�z�WM��d�A�k��A:�t�+⃓��� p%�:���5�]�S��lg������!�B_��{�FZ�ԕah85͗���ZP��d�)��0�������ؼ7�e�L߼��
�d{�<P��u�D�
BJ�!ٟ�Lv
�<�?"~�E]0i����Ѩ��?���S��/��T��V	>u-V�o^�<��X�OTO ����`���6..�q�B7/2x@�����L����ǷK3|[�oB� !D�����x��n�A�N1@����p��i��t�+]�'.<�qYЃ����D�<%KYn�n`=W,�48M��؆_֢��O8O���b�4G`�)y9$v��{.��d�Q�(~l���sۭ���Z��7A\��v��]3��#ҩ�{��)�vA4�F���D!�}��I����B����m��5�6Qg)fy��fR/R��3�nt��tzu�L!w9O��Q�]گm"����!-�<޹��Y"��b�.�)�nW�!b��K4z")8T�2�f�b��������]VJ9B0�����Ƹ�������"�~b5Wg��N��sH6zU�s�_��RG8���q�F�XlxVHYEB    9732    14d0���M[�2j��ˊ���OkB��>���*��`�j&�������N��V3��h�yn9E�i��Q��|8��f�//�GST����$�!�A�~F���J���X�ӎ٨9�ir�y
.�c�����T^Qu�6>s�S�:㵣S��L��!���a�n�-'B��ON��C�Zc��W���{�Ä�HF���t@��!뫏L��B��p7��
���C�v��3�!�w*	��Z�����2���=J

�8�B�,\F�C��8�Fќ�V=�q�C7J�V:� �繍�}�r8c�G��.�&)�tIQt�\.����'�>[k�dY��%dN�V���g��`.����P��c<�3�\c;}�B�SCD�~�A�u{���C��3C��\�8�����f�W�?�&��%��ƈ��k�w�m"�ɸ�NZ��ܴ]s�����W (rł�V�r�6�Ț�P�!�\�/���p�7��&~��ݬ�K�r�-���Za�;,ݬ<����*���B��8�r�G�j����	Ҍ��Q��о'��sj4����H�V�Q�*F�"a�����S4J�]�H6�{$J��Rg6�a���(��Jˇ����8�@�͟f��c_E�����%w>����\'��9��{��l�5I0�G��J)��Ѵ��'�#C�l��k�!ǈzc�b$�2��8����[X�y}���_EQ��/vvB_wʶg�?��ӧw�����[����7��U&%
 Կ[忬}��e��hGbLs}3S.�Km�~>l(��x�W��uK��5~ʁ5�Q�fS�Uh���oڠ�W�h=L���'PQߝA/~���F���������1{��c5�PF@Z�_?�)�HV9���Yg��A2F�F�0�9�G}��;��|�TZ�Y�\��R�i��-��@�����&&MC
{iM�S����E����QM�p0���	��H&h�jez���nӦ�,R��Y�5iR,@����R���ݎձ�t���7�X�S�v��+�(ί�ZWCR�_�BS�[��c��3�����t�l�r���`���W %|�/���E��V���ɱC��b��y2@F�P��=D����&�8|m���s�r�<��k���������<��'�L��
x$v��~+#�k '�De������U�H�-���Zk�\x�;P��7!�%�3]�@AK����
�S�VҶ	���]��hb�߿:շ�Äɐy���g��-�� ~�[���^07�����(�B�8��X�!@ƺ�V���:�X��ʙ@w������ޣ�`V�:m;�q#�Ǉ[�h0=g���9�a�L"4� �_�R��\t�!Tʐ#R�!N��ƫnEPNe%�h��AS�y<��L���k�4�a �A����yF��5W�'�]~�1U#$�I��3PF 1�j�1�UP��-��BRP�"|9�K>P�JS�Hi	���U���	���;g6�9X!p^ƸL�A7WtӀ]�Su��Xn��h#���H�|�D=�ƙ�u8C��4��=��K�W2��Kܡ<ni\�<��)r<�N�ʮ���J����жa��lL���B�/eِ����N��8uT�5�R��������Yx8O('2�p��T6en�0���Amj�Lw����`���;W:_|�wZq��o��p
�Q3��9Ҝ%-�Rn�<7�X���v�M��S�/�� �=� ��Pp�p���ߜ�ve'�o뤤$l��5\�ֆ���s���g$e瓜�[=n�x���	I���䥼>>�
�[՘�+�nj+4�H��N[�q�pd�ȲX���:�᠝������3��zԄ�h:w�}r`@e��ݏ ǜo�����Ϡ#��O��-�"��TC楮��9tƶtC�E���)Ԩ�H���O�^3���7�o�~��~������
�l���
��)l?� 	��FZ7j��Ƚ��	�QcR�^'�U�L�3Wc��
�"C��ͫ)�!�<�%���9b��g��`��J�(������ Ҡ�2�|#�9휉�׈JC�$�$|��w�&�82w������e�sF��mvE�P����{��]g�ɖ�p4}ٖ�#�]a�&w�L��ڲ����oɜ~��;zi���~H���뫏v��Ǳ�)����m��^N7����T������ʱ��[*�`�-^֔e	O�-9f$��=�ƠD�D��V�kv���M{>���8T-��4��ߗ�K��חq#Jm�@�t@ ,˟C�M�SdRG���%�O��:��OƩ��̳��{ԇ�V�c,�]�U��H��ޟO���q$VSu[Y��j��Nݟ%��g�����B&�_���3�������(�#EU�Gk��޹��7%��!��|`�[<J�Y.���h
Ɇ3�����D-B��!��T?���5Z����O�J:��U������P�`4�;�^��x+'je�ľ�A�~|%��>�:P2�w C��&�*lnI�����{�[�[��{��R���[�י��ʍj��l^�Ơ��I�B����>8�X�zۥ
�=qY�p{f��[�>[l!|��G�(g7v�S����¥8�ٌd"U٤y�/Tw��ƌ�t�*b�x�U�)��?ň�ϛ"UGsrgl�Se�$v�φK
R�[kO1_��k18&^p��x��y��Mr�F��v<���!_A/%�L�L��h��:���nW�Yh��5<T�}$�9K�����QK�`�<���;\Rĝ�r��H��b3�"y��:oaI�@{��cc�k��sz���Ge���%\�+������辀 Sl9R���t�8��ȷ�5@�  !����G5ˡ9�&����l,R�'��1��ү�d�X���\�$�q5����=�Y���Ɔy/��bGc�ɝ0��̎�WLR��_��JyIO�\�����y���U�ٍ(������Ј�Q����'9tMV#�{��|~ɛ[k<����oK���Im�Wo_�̓K��i����G��ŀ2#���[I��Vͬ�2���&�'��Ę՗�u|	=��*�uQ]P>&՗.�wb>
0�N�Τ��X0-Q��(�~4�NWU��Ui�6�	���+��ƙ�ނ���d=�oi ��c7"/6O��A<���^�%��T�� ��M�Gv�2����D�^��ⓜ.QG��f1�7������K�ߨ�i3ZSYY�=!��E���RQih� �<ȳIo^PO(�UI5���j������,m5�/r؁ ��&�%P�h�/�֑�)��5S�E�I0_�ԁ/��4S�Q M�]FC^���E��u�PG���4�hƱ�-�H�t�#*���QhFTRud��\���i��?���'�Oet>�(��{��Ň[)�E"��k߲��&���'���i��F�Ы���>+�"`).����3�!���������</Ou�������|�L���z��OZ(��
Ӣh|Lꇬ9+�od���[<�M�X��f'x�s�h�������G���#]�t3��Ga��� rݫ�A���J�K"mt*`y�����N��L52�ם�[i��J53�����4��!�5��C�t���eߚ���;�{�$������W| X�Rn2?������lc�#Ϋ��}j�6Ij�I�8���_&�X�0��l]m�w�і"�t�T��1��e�m<_�Т!M���iH�}��8a����j����#�&����>�౴��w:8�1m7����M��ZY�����˾M�-���s��a�#��t��T%�?�;���Ȏ�q��n���L a��n�¸-Ǐ}�ΔlO�Ֆ����N
?�{�q��G�첸W��I4�#�ۛ浴ռ��J.���i����El�ȈS%�^6��	�ب�|k��㵘�k���%وI�y��տ8�P��z�e/���b%M󣁔��Jk�7Ց��V#.[���y�K�k~=9�(�Ϩ�a�P��@�{e�m��T�?�n6E�i��Lu��c+�`�<a�ʕ#��de�L��F���a�>�u�/�v�Y_�M�<�hC�qZcZ���Uߋ��s^3nr/��i"!K����t<�/���l��6?�w:,��
�;?3�D�>�c2X Q
�)�vخ썶�
P��l�Y��54��g����w�=��O��i9U�c�醷<Y��G��D�o�N%^���g4ڻM��w�Xf�W��,ױ�B���#Mf`�đ��z���	��
��T>z6d�E����w�#3��.�&)�I"5#tً��$�Ψ����e�6�/R�H1w+���ho>��:��	F�ڵ��oL�8���m.K�l�*~����uU��� b/O�� �ÄM��]*�o&��,�Z��u��q�.��������qr
��tF��Z���"��Ѵ��
�cr����B��c���]~��Ƚ�Uҹ�'��oЗӹ�ǔ���?o�
f�(�.;(с�.��/��e�z`���v0r��)�J)x
/X���O�ƌщ�k�4;6O��3�����U��i������sA��� ������k'�;X�!
j��)��.G�{ �[�8��W"��H�������q��^�n�1;A�rٚs���X E�?A�V�g*5� ���؍<c8���}& {�a/��z	V�+��^���Q�a�ُf;���BN;��pi���i�zf��?|l�?-��qZn�R
�u`����b��
���-�"m�����|�[��}�b�ZI{�@ ŅҤ��ƥ@I��v�B��w�E=e�h�V�Q�Θ��$H���B�+^\h��<a��U �l��mqG�>�`V�E�Hpon��9�h���I�k��Pg\uHW�6E�+�J�yJ���<h�.����qf�"�S�G+�d��le�j�8Am�fO'0l2 J��b�lI�NA�����4'FE$�!��[sֶ"v.�`8s`%�Fpٙ����Ro�jݏ�e�c�p��04�Iq&�c��D��t3�F"u��|��Aү�\x"jݖ����*o�3�Xx��4Z��ұVDz`?�3J�܁�t�Ց��?1-��`ަP,1�B99�a��~��Ї��ll�W�׷����;8�O��9,�s7��:'[��}Q�[�9"G�-�����S�H�}c워�v	hi�����
���C��*Xz	�ld/��ֿ��E0�6��^w�����M����/+�t!�I]�ɷ*�NAo�!�Q�6���>!���$�)�۰��n �.Πu�8�	�0��V�~T�r#�7/��0��|̛�ja����@űܒ��I]�嗿