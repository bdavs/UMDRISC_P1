XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��FA^�#e��r`�q8u	j#�M����;/?oVv��S5t�<F����,8�ol��|cX��~?�9����?0"U@'��\�PqJ/��W�mv�t�,d�B6���2P�C����ƶI ��"ַ����K���eP����r��Y%{?�9y���]���e��c"J��  �_�q��98/&8�5��s;z �0$Tp�����`M�E��EՃ���8�ڱq����Ѻ�
}�ͱUQ�@������͓����%����ס�v��تO;���+�t��D�[qC��e]5���R-<Ǭ2X��TA��#�,�]����X��"�����t0"=��Ǧ`�;�C�!�>r&ڠ�vR��?aQ������u����-���7ǀ��9`�2�^���
������ ��;�J�\:��4�	�%a�z�V~B�d"�q���"��9��)�~�#^VL�|�v�T)i��K��r�x�2ĩ�P�e��<���x>��r9aTe+رF�{�Z
�ԙ��p�Z ��b���!��%��L��L��Zl���e�#�� �6�SȚ3t�%M2�`A�b�b���ZۙG�X����Rw�
IT��ȅepS�L����18lI���2������bt���{�A'<��m$���\���Oa���<�;)>��K�,����k.kW^S�!�?zW��7`����6����o0ma����VF8�i�q�c�n	D<��� RزG�91�y� �d��稞��b��XlxVHYEB    fa00    2950�{"��l���|��aK<�ʀ�fk�Ƅ�������F��P8u�?o:�H�(6�cMS�@MpCS�l�rlt
':K�3���U�:���v&�,�Ḥ��ҥ���%d]��O"ΐ��FT,1��n�r��a��O��A���0~�9���f���,� &�u��y0��1��抌N�;D����SJv@�T_W�ή���g���'[�F�a�ld��d�C�V.�B<E�3k6�[³�ྤ�-�I_�Z�w��t����+��},2q0���l��ed]�.��y�V�w��u��_Pd�J}b�BP�8��n���>�Y*nrӸX�u|���q����5���� u�b����t��/�Ǧ�^���B����k�y�%f��Op{�^�N�Z9�峃q�{���� #��<�F,�{�C?]qAp��H���������#P�7>���Q4�̣�({�xܧU��ɨ�̓O�˶x�JT�h$k5�[����(Y%?w,�P�e�+w��B���=�'|�A���ј��/Ă�]97��a >ށt��j4�����-� J���ݶd��5\���Õ��Jx�V
c"^�k�hݻ^��`���殂I�k�H:��@�^�ķ�o��UG���9�Ǐ16�T���P�C_@�t'F���pN��*��#(Π]�����6�A�SI�~�K�5�g���l�r��Q0���J� �u��@��b�IHa͛�� 1Ĺ�J�![.q�ʻ֧�Y%˳�+�@`I���N�J��Sۓd�Xk�R��P���fʫO��v�mbQk]P�+f)�Ԑ�ZO��I>�Yl��/���(҈`)q�An��u�g��G*�M��$'�6F�XU6�ˠ��N����(���g0!�ś��Ғ�n��7P�N΀ߊX0�H��d��)U��8�U�����o�|,!,۵��>��I;�/�J�����s�����I�U(]3���6��i����5���G�ix�'�x��/�'� N�/�,_���p���f�~����|$��/�^_0{�s��K]��H���L��=�^�Wk5I'��
Ʀ�l,�_S�.��Y3� �g�Ez�4ǘ	��hu�=E���Q㘞�D�(� װ�D���
��nr�"�7��69~���0�cC�8SS��k�O	���Ъ#���"G}/)XD���0}���i�2�妑�sI���1�U��ݏ���Y�t��T`#�=�;ٞ�N�����}�x»	+V$RZ\�xD|����-VH�R/��fs�X��8W��;Y%�9S/�;�P(M���[��j'L�O��Z����>[�����F��bdO=�Fh�#a�k�:�#t��̄`y'i�����ozHC��jiF#lSi��߸��p�`�|E+P��۱5���2&Y�ꌸ�ȶPK�����
���m�AE��?m��4��$eF��ɗ����	��A�����Oj�=�0�N�H"Q`�-#s_���� �t�x5�����jN����掿��R���}�o���G�X�BFS�'�� z�Yv	��g�vZ��n��m�s��^wAM�t��W� N-˻�t�A�`�{����-�w���}�{�^��6�,J<ۧ<�߆�x�|�@����PY�Lk�=�r���|>���|Eٯ�Î֩�Ex�(�8�%&},g�f����
rG�&���YJ�J9��SQp�"�&Î2掟l&�w�_�4�ʶ���yM���M�R���> `�����$'��O��
|(e���˹�p��cΐ@�>�o�*B�2�s!��j�YS�czaT@RI&�B��:��];��ct��Q�j�&�[.�7��3f�88���4W��yΩtG<.9��\��d��΄`F5<j!L���~�P�1����Gм(�J�kV�})�u�O>2�Ǝa�%k~����(R��pO�L� ��H٠�3��N5�P��z�����p�wIS�q*��46wQ)
.��%g젎-/����W0��%�xV����_5�Y����􁥣`����f��C2�^J`oݗ@�d$��;$7���ؓ0N��Q�N�3��'d�^V�s��n����r]-K���T,��T�����w�M�9��M���*j��6�*�ds 1�g��`���.�6�.p�dd�?�	&<NW\�����+ii�u���;�Q�Y������w����7�Ӗl)�5�e�:N�U�PN6x\�'���	X���Ѥ�5;YB�h�Oqa��
�Q�v2��^[������I(]�Z�$��~�%j��A�R3�N�塚�aY}��:�\u��d԰p[���u'�]|���$ב�4�)��r�\��Nd��CθZ�q��,��c.'�"���_[����%&,o�TQmJo��xR���L6q��a��Z[mT7Q ����|pvDo'�һ+eŀS�p�.-Õ���vo�칑����$°�o(�c��Q*\6�9�@�Պ&����RK-Z"L��{9����s�Xͷ�<�{ya�p%�(������'P�>���/i��@T�3|lL�TG�/&6%���	Ea`0y^����q~>A�[㽲�U	�Փ� }�� @�s�na�uЦba�ܺ�
����FL��ҫ�]'8E��D['���z���i
��W�����M:��tm�L��2K����eh����I�i&ʁn�o����7b�ӟ�[�jL���j�B�NN<�8i�j��ub����>�Q������a���~�Ԉ���l�n�&��h ��<�@ s��L�D�+|��D+��e�n�hX$^����77�Q��?両���Щ�أg� ��{p�)}��m�v�4�0߽)��j2����Xi�$��i�N�ܐ�~�'f}u���,�j(.u@��R��k�{�S�5�5jW����M�	c��E��G(�ђ-:�f}��~sEQ'�KsW��U�/�T�3{=��\�"f�[f9.�|�U�*��r���� �� xA��t_9E2�D�AGW��$�
�����,ޚ@� ��@އ�������q�< �L�6��P/w�.Ӕ�]�_�IM��	��\�$�"��U�L����5��e���z��[��.�����=��(JaJ8Ȗ����?:J�������19`b��P�E}�+��������b5{�a�I��?�,�7���I�by]��׮� s�5��M���b�A�f�T��ځ�~vB!q�S�T�(���ZZ�`W�u�>�~�ڶ�=�O�!�,��B�3���uFb�-CRN��.c#�	�ίpiGȮ"R^dd�Ă� E��W�!d��8�4�<q�QH�j�
k,U��ӫRd�i%|�Z&$�O�LW�k��I6IK��cF��.TO���vX�h�v�9<"�ܗ�6"3׮�T�j>�h[��!q��&������]�Y�/Vޅ� 3+�;��+�T�M$�3u���!Č���9|i�D(F��s�<pbI��� �I�5^$^���
����dDHY��⊃v%+MG�sM��X�?�خ�����l�t��Z ����Q�P���]����	ϛ����-Ts��,�kF�v`���H>� yf�gf��
�� �a�_��}_�y���-��o�`��)I�(QߺЗE�iЃ�%0���{;^�e5�  F�i}�B{�MWz|�'U��	H�����6W�Ttqu��k�c�Lχ�e���6�^U����^O�p��$\�}\j:h;����V	;�5����M|�nv�٢3z�{?���?��Y�������� ����(nmM3�N([�=�� ��T�w���-y��x�vS�2	�yn�DDS�� �(7T�!g�%Z��J�/E1*��L��������e�Y�.Z?���AyՁ����%l�d/�MЦ\��줍w1�����(�$��e�͹f8�ZD	(� ������3�i�pt��ޣ�@l�/ba�-�S6OR_+��ч����z��~7�����A;$�e��&��7`�+"ڒ�X�% uy����l�j�i[,�����"j�b@P�g���<��(%�^����"�7GxZr��T�P�(��&��P��9E״$H��F��~��+�np+������6�0�Y��=��J+s�0'��8��bB�D���1�
M�<���2o�J�2_� �/�em�}
\�������f�Ci�h;�yJʜ�CFP@���Qv�&{!ش���7,OSbd�r̛_;�W˽�E���8�7\��_i�H�`4$���0r�T	�`����K����8��Nm:�!��qV.�r�U��eqQ�n{��vÓ��ׄ�b�����-������D+	���=�K��M��kӍ�����ó�zE�(�J,i�y�l�X�*N+�'���=rd;��+D����ލw3�q.Xʵ+[��6���B��+۽���[����) wd�����&�7���	 ���6�Gmli(���g~��ւ�n5����/������"�݉����V���1Ly��aE�Iζ�C�(���X�zms~r�܋��}��� k�P���6�H�JJͱ������]�2'G������ҟKɂ�����,�M�@���V�}Ai�.�V��JPC�4^h��'�080Z��&0p��p"a�g`�,e�ة�0�>c��{	�Huc���������oW<�1si��-
�:tF�?���[�&�atj��8�.o���1q�/�	�$@�(����tWǆGM���Ԑ>��ju-�FY�S� ֵ}"�=A�#��1��s�ї�]^�?��IgY�f�3#�qÿ<._
N����ʌ��(?�*Yj�L�/2d�sE֣;\��n�p��b��n�O�G]�J_�����G�Q胔G�� [!Yc��U�IoY�;�*G4a8#��|�)Y���ZO)4�"2?W~�ͫ�Z�k�m����5q���P��V��2b�4Z����>;����ٲR׶�|N�/=F�}�h�F�h�������x���5��v���_I�C$]0�ֈU�g꒘H��$+!M<��zT��N�~H��i��?����	-7m��A��� �O&*������S�ؓ	�Xo�0;^�����'�B s��;��ٱ!�:VW�k��*���� {O��7FlU}��h����Lq��[]Y���ZU��{�����_5zJE7���lh۵�	�8��!��d�H����/K6�"C���Uo�"�E�U��L��h�g3���YM{Ԋv�r7�,Ot������������·j"�Ft�������M=B��laRd]#>������i9wU�s��Ũ����ʮ���x��W���=��Tn�2��ߏ��a�_���\��c���(� ���!�v^*�줓��[m|��`f��JpAK���%J"�6��fx�s�����m�A`���/$�[	�|"�F��ah�Fxђʸ���%���:�GJ����*��ՙ��P~5r�pA��I��O��G�z��:����)W�,Z{T���1s�LX<1��u&^��s�]m-��T�إ�/�0bCd̐d��^��2�Kn�$�H X54|����Rk��Z�9�@�ȶ�����VRO_�2�ơxB�Nm�U.o*?�8��	#��4{y����\3���g�i�|f�4J(�������S�X�J�����������}S�@c$½b�m�ye�[�.�T��y(`��Oņ9�����
�[K`8����f ��|яN]i�防@/������C�ب !�<��#S|�{�,Mc|���.�\���'|�HNj_p8:@|-�����T�{j���K6�ҵ���i��m[Q�-PLH��y+Ba�0|DF����zy L?WU�{3��C�h�gV��;qCEG6�T�\��s�2'ǔqN����7�y���!�=f�O�9�m�
+?��IKB���n��^��XH"����:m�����1e��O�(�6C�A����\c�aG�>}[�`�"��m@رRx4Y]G��F�(u�|�2n�K�ʙ�(�K0\�	4K/'���4��8�\�I�K������R�,M �F/Y��{g�C�����>z�y�� ��˔-���Χ���.V�Ԍ�]n1I�,06L�j14��WRh���@b�{Q]��*1����$���4����]w|ߊ��}��y��ހz�S�C�D��r�X��*�����'���s~�w1�T�k��>�>��Z"�e�M
�j�+�E?�V8J�_�}�U���;־���깂! G�"K�[)�P�j�/G�&��(M�?�0�F�P{�R�l�	"ty�րi�U��yS$�_��}����0�v��	������d��h��|�3��)9��?)�8k�b%B�_��=}�}���Dv�Y�(���I���`�Q9�aSG��T�����1��M"c�%	!��5m ���y1�CKR��d%j��a���V�#� *J����PT�,x}�8�Y�K{C����H��*�c�P�Z�wF{�-)Jd�MjU����GH�eU�>C�e�L)-� ��Bˋ�>�%^	��������V����3���;`.s����	V�V*HZ?��UFg!.���yN�U�����)�ѣ;ֱ������0��M�.h��G���7axw.��]��3�@���Kx���̳$KT�@��U�����P����ŉ�/։�WZ����'�"��KA�m���8���3���n�>ڇ�ӹdr��~[3���Mh3�%�Pp�'6;(Ծ�!e�zM���8�bv�
�zz^��J��F8L������	ri��&\�L?xUc�~5[��p�.�爾#�@kŞ���مm �H_p����G =ak.�AF��؇W� ��ѱ��~Â�/�oY�3��BtJȶ�a]�kl)��&��l����'}�뒫�'eÜ�U�D�,vy���;z+oY�ֹ3�\OW^��S� !V�"�����y�����No j%�C)�����~=Y�tF�J�(��N'�"�����^}��:�R1�5�pWh2W	���P-&�����,�F~M?�6��pl��b�8g�Y.dȍ���~���-�z}�}񢋪���?킵r^�>!m�y/;8��s��#ש:�U�w\=��g4>��	�������H�y��A�h�{�����<*�Yg�d�Ɲ��d����H!P��p�X-����.W����1�7�����&��� i��2���H0o|?�rѩLi&Da�(݃���l��y�؍N�J����I�:>���Kf��E����8S��\�o�$����W��P���mK�ˋ��g���g(���:X38�\n�5�]�&qm�'V��E"�A�#[��i����9�ॆ{J��xwM'���R�P�3n �5.��ͺY�Xކ`�еVp$�&
�X�ȱ,��Z�tQ�M%�&��!N�Qt�֨��М��ey�i�&ܑx��r��p�p� m�h8F!�R�G��g�>B�U^?w�`���?�,s�8qY5�rc��F�(��~^�`���IV�~U9+4�/�v�����D��R��vXz�$_O�EQ�m��2�q2�$K���Ow(i��T�n9��n~#��Ux���xF.6�}�*�8}`o�6���zlZ���}�X���h_'����`�����05ݐ��y2R��=X7:]� Ǩ�����H�(���P��C��c$O�#t��m�#6�=$�&L_W:l��H�?$���=��QK��<�~e�j���+�yCZv�R�)rXa��/�X#`e����h��f������n�a̬�k��D�OMg�S�J]������/0�^�bK�/$����֛��f23n{LT�D �W����7��ҫ�E��&��P�/˷f��<�M�c����k�.v*@�2�>X�D�.��d0�bʮ����Y|��0*z�;J<��5����u�ʴ�t^P�l[t��sZ[�j�f�oڌ?T�<�)�Y�Q�)���C>zv��w��x��SS\�}�I�%����Cf1�D���Aw��CA��|��_�0����1xY�\��;���Z�fчm3�b[�?��0(�� ;�δ4A&�R���4i~j���{z���+N	�����&�ŀ� F�$R4S+�D���*�P�*Qu��Ԇ���YK X��v0�Q�דbG7t������e�])c��x����eI�0�r�M�k��[�e` �0hf�n?<P�׳;�cOm�)QY��g�uHF�������v��g�/.�h�^1��[>�" �-q�]�E)��-]���?E�3�-����%ѓ7���3�^x;��GCp��^�k|;��4���r�(�Pl���9�Oy��^i�� ���LV��M��i�n� W��i]����b4)//i�ښP��T��ա�;��'RGK�+C�
�S�*Df���ԋ��Dx��3=���Fh0�D��t����6*���f/%�,�5���le	��sf��d�hpug��֛a'rSݲ�{��畐����+�Y���0p�,n�����0'���)�pɌ���e��~y3H9�������|��w����>�%S��و��Gk��/�z�<J,�3���dz�A&��qS�����jQ��脥=b�cjr�3ʕL�+�jٞ��-��$�E�W��-F�[ŵ�L"p��s��Z���z�{0/�,
�{H��ʄ����i����V�ʃ�OJK���Zka�����a_�$�h������_Ƙ��KZ��\e���W_�/�Uj���ʊL#<�U��@��m���A�K���R��T�0B�J�_>EGh0BR~���)�o�((.z�#�_+�2)����Yo�A��`�^7�����|(�j�c������Z�z|ZR�h���v�烣\��p��8��Z���t���/�nӹ��ð�zT	{F�'��r	�i	<6ն4��������+� s���b��7�^��(Q�z9	�Ef.:�Bz!3]�N�Qm�q�a���K�"��7gZ���;[�ks�п���K7��5}���������^�yٳ���dUFTLq����ge��vtj
�k�TV� d?���4�`+�˨X����x�,�`��c���}=fH�baǳ
vMd={�s�K�"��R�	������9�]��;��A���Km	�SېΡ��(��k�&��aC���!kV�S��'�ϾN���)�% '�P�,�|�O��>7p�g�;�	�85�UpK�'_�����˙�jsZ:��S�s[���}�m\ko�3d$��n��>��yMpcݔ0s~�o5�<��j���A�6vAƣ����p�?J&"�v�쫦�e	�!+���D�AY�	��ME�y}���p[ae3$z/D�O	i�����V҄��0���������6���i�����&C����J�e����L7S�4V�:SO_�0��}g"3�a�ʴ�}�O�C,��/�$�|	I��Ӂ�Y�ܙ��:WAW�In�(��`�qԈ�H.�K�SAC�y��CW�K��~���U�p������5?���U��A����,�$r)ܟ���?]���T$>m�pʯ���yo���%�a�[#ge�CL�B�*@�SDW�eL��Y�?L�Q���A�?f.�o8�s�7*�i�gwĺ��`�$B�v2%fu�x�:�a�a�
R��ş��QPdWDj�sDH�L��#h�v��U;/'ʫ��+�Q�Lݟ=I�e��ԥ�چ?o7$��������z �&�/�5��^����+mD��V�J㥉s_؂���uS�"���Ї���"�%����+r��������e�M�o僆��(�$���O��5u���l
���l��D�8֑h��.���2u9�Z+��d)^=`E��sm�Y�*m54[�	e9�f^�k�}��W�\rG)�#n;�Ƚe^a��6������S�wyv�9�6l;��y�	~����!��`��"��������fKJ�D��\��o9�2pz@;�m����n�
���գ�z���-hj��k�=�/���0��Y����ӌ�xc@�0g�d���A#�K[�C ��
ϱ�#�66�R��s�x��4�:���Ep�(� H(,}A҅�Z�I��5
*@�C �� ��z�Kܭ�ӝ��P�v�������_�i��}��<�3lO��}*`�'z~hQ�!>6v�8��#�m8�����_�O��I�S�9���k�Ȳ�t56k+U��E��8Љ�Ȳ��*� ��z�M��g��:%k���p��g�[�h=����r��$�O���_;��4��z���1ʺ}��S�0�es�>��=
y}��c!YYVlh�T%tgZ2���gޢ��9��XlxVHYEB    fa00    1e30lGC�:ι
�4ӆK�񐿕?��tS�j��a�D���F��3��*FKS�.�����=A�R�I�5s��nȆ��Y!�>��>�1�l�2���Wi;���}[ʔxX+�8�V����H޼�[e�`��~
50U�iH�L��&SDMVw1�q򌫠=s:�]ò��;���ܙrx���ѧFv{�A�
}�LN\<Z*���$9ў*���8�|�a�Mv`��cZi��ok����Ǹ|e�dAZ�d��IՄ<��z��Z���6ܵ�1�o�������q㻢F����_A�3H�������@�1J��C
�.�8Aʰ��;К�G>9zg��<������w���_���Ӏ�g�x��lh}�y�}w,T�qKH����LI@�Q䲮z(��5�����9wG�hS��Qe,H�0E�8��cw��������VR$�Ĩ�\>NYϏ+���Gr5�0�O6�^�L6��:w}fMҺ�¥5iw;f�b�0wg��ǏCܬ���"8yUF�P��F��3	����p~���Mg�)��4�4�[�_���>x��;X<����S&�;-
^����J�\�a�jW]3�mUMj�RMĞ�5��4�Y�#3���L���ԅ�h@�T�*��;'\�?�^\�(�d�	ʽ̕�W��_Y��N���u�����X���q��ާ^��'?)w��p��/|%�����(!h����C��:2���|dS>U��d%���FTPb�?��"��g�*��)%�_PA0��x���=��$���7M:rG,^�C _V��A�.ρa��u6(�{s��G��iq��D�׊��x��+�kt��n���}�X8K�s��fCf�J�i8�9��U�ݴ�E�컫�0���F:o�{et'��:�������m$��HT����Z�^����"��EJ�y�4�Zm�_]tb�0��gp�U�?�.��r�lT&|V�%ўK��\��y"��9QX�@���^"Pg5]����C˽=�;顂+����X�� ����
��2�\��ɻh�1<��SC�֑D���[ޣ��!A~�*��`�>�B�ҧ�!�9kuT ̼i.�e�!���R8�ѕJ�df����c�z:��K[+�C��j�x_��.b��L麚b��ܶ�����D�#�ع�b`͐H�bC{�Ђ/�VT��`�r�����Up��t���pw^M�<[��`�����6��?��I��������r�:MK�XD.R��0n�%��ۢ_iiyM�L�\vͨ'v���*��3"��?��r�;m���.z��6�ȯ���=��v����>x��xɠ/�o�+M��1�B����PUA�U����b��FW���y���-"��,&�����T�Va�P��k0:>��B�)`@̷��,e)�&�rD�b^�U��kV���
��	+6�n�?l��Lٚ�'j�C^���������|J����Բ����A�ě���{��9zp;�N�.#��)f}*���%�~"C�/]�M�V��2Pt+�Gi�%u���#ߥ�O_��P-݊{.�3hy��ʟXhe�h��h2�ը�C���v������5Z`l�^S2�osN:Ӥ�(Y�����j�l�ㆀЇ��Xv�_  �v����I�В#]p`�܅t9R�Iۀ�O�ݥ3V̀bZ>� �NW8��3S^q�[�;n��
-Z�F΢�1�V�	�:�N9A��t�[�w�S�6�#Z�+������s�����1p�"�<R�.H!�2�v
��I�R7y[���Y�r�Cڶ�/1�S��	��InƮ
+T�U��s÷��<Z�A���7蚓V�\�M�������M~R�����(y��(}��'n~Z��B��#�ڐ��������F���n���c*��G�N�������d��`�SG iC��a����3Y �&��������/<V���0Խ�����2�ȡ�XA��Tt@���O��BA6��r�ߴ�⺳�j�/ϣ�B�Ap��2�[n?�2�y�E�ҹL�?���W}s@$�R�w�X��I�O�1zs�ϥ&���bO�;��MӰ���׳��'��8v��^�߾���>��q`	�O	Z�E@���F��B�&���8���=��l$e�mg�N��L��`���g�5�C�ty��-��Sf���ik��o��M��/��!�����N�i�,��<�BN�P�����v��Y���eZ��̙fjXy�%L7����/ �Ȫњ�G��;Q�������:Wƌ��/�ik냤�<�M#��������С�ia�c��O�3:$C�fh�S�5��y��<��|E�N|R=�PZ	aPD�h�����E��ny�T-w��Zqd6��/�y�D�E�Z� �}��eA�a+}��0��3���Bc��z`G�Iq�x4Uk�����U&�Qa4�O)�	7hWt��uX��*�����:c��n����b߼�r�">MH����mI������G��Ż�,53O��BhL�g���_|G��Gj��=�#�"����@G<{��gh�*����2�{?m�b�-z��R��|E7��P��
��B�=���AB�W9;����%�����7���	΢�>�ޛ�d�����u���lw���	[�Z����+����>�!���(Md�K��['�g"6kS����x�O^WX��"�.oߍW�y�>TZ�G������
g�A�Y�*�FJ�F�e��@)��.q�^��[��1By�+Հ^��w2G#FqP��ͫ���
K�Ղo#�tI�1B���y�u&�37��v�zx�"��ϐ���N�%��;��0*Q (��6�d���?����zw�Hm ���@�� ��e�V��P�Vp�GH^PXK>�A��#۷��Q�|�v��T%�E����i���A��� ��$wp݊ �j�$�y�����'��N����l�s��Ԃݳ�F�>�nM�}�Yi�+��ٓ��	3![����3��ʄB.�@2�HP�M5z��ͧ�����hZ�Ʒ��	��X<�벷X1�"����mU��6;'DP}�=6�Dٴ`���6��a���ñݿ��k�B$wK5dM�鞕f'�UN��,�,�X�gPA^@�s��,[��뷏��s>�־��YϮ�n�d���� �K��;��Z�����os�dg�Њ�Y�RC[�ʪ�i�Л��߯� ��EV��a828�[<��k��)Q��N}%k����xH�6V �~�JZ�=�F3��JC#(�!�MS�=V����}c�������|��r��*��Q��@��Y�� �J����n�jf	'�h}�-v���?��"��|E�A�Z���#	>y�M�	( ��-�1��Y�Cp�dml�#�oD��RiN^J�������F`�:��u�	�F��٥���oK ����_g~�ؿ�|�\�/�_0�Q���<���Hh��ט���pb�N��i��a��+���[Cv/��0_���3�1�[L}w���_A�T���gbt%����+��{������^L�v�
h��N^*�:e���}8�K��VR�tM#��>!V��6x��v�	�6�/��!%��t%��h
(�GW)=�'���K� �< �n���&��{M�"ZҼ����@�T����H������sӵ�Q����FBfm��
���aܸͳ��|�m{�=�� R��!/ؤ���6�m�*��^��d�6�Uc�hJ*[�z�WR�!�h_��R��E|��TpL|7�˶-�@��*�;���cz���B���~�f�H=.�<�
*�M�$�IoG�~�fVxYTb �ȶ�Q;{���@�̗i�
N�,�L�� 	#������C�Uu~(Ç�b���uzur�Mj�N� Ի|ƻ��_�����oX�Vf�N'�����m?\ ���A߹?k3�8ob&��r���f�(a؄Eso\�g��t����h�^P㛢����5ͣ�V��3H�H<b�_S�DwCI��d/�2^f%�>ZĆ���y��ا��p"=�GG�m��w��Z�G7��������fR��iPK$蓫K,@��HR��މ*@���8�=Bc��|�gX4��_n�I"���4���hjᎰ� ��-���l�H�n�������(��`�X/�h��,����ܱGE;z���=��׳��{�ϙ������z��@fט����x���h�7[G9�o��Ǘ��k?��|��'}�1c����Qe�E#����X�v؏=n���N@w�p����4��Q��,�����C,'���^F�q$��>(��a^A�6��h��{Gʍ� ����ӄ�O������<,0����~͒{3L������/ߢ�����_\ښ��§�d�HaT��k���Ӭ���9C{�����
3x��:y�����u>	��?/�o�2��  ���%��p�jgS���Ӱ�rb���v�O�����wq��߂��Z&B<�ˣ�8����NJ�I0�U�&`�1�T[�N����C�ћԁ�(�e�`.���H	�o����?l���Ӭ�9��^-�5��r�36iа�k�
�bJ���#�E/a�B&cɛ5�S��v�J�zym�&ǐ���pֶ
��O.8W��wO��GZ~���-�B�9�S<[SeA����"%��H�vǤ�1��b��p��q$ ��<�)}A�G�B_h�ImE��l���y�K��릓�,�D����:T��.M�wO�	vN�;&���|`��W�ש)M/�{������#�r�y-��O�Um���(-��I��a��9��%��l��e;�6^�,$��C�9@�2��X�����+8��N�/޿޴GE��߫s�`��܄���E�]�x��^Gk��ex	�_^�xyCh��x Y'ߋX��d)y�<�2*b�������c&p�b���D]�w����K�� Iy����YLlV��K������P#��7�f�������)�7f.o�����b����,�V���9�
.�~VYA�ћ�ftk�l
��0 �Fy�?-*2�O�)�|4������^��g@�`�qz�S!(>��.�ފ��~���X�����X�*����&n�Yo��� ,{;��Q��n�ܕ���䑯I�-N@��x�f�L�%�Sz��p�$��m��qˇ�G��!9�B:����\Hsx������������Z�CA�-�:�-N?T��)��c����ϪOTwIh��z�ēt�Xg��v�7�X�0^qS>���{
T����H\��5p*��5�����=|
�σi��G�����S�x��6j��R�$ϱб�LV��=���x�c�����L~X��x�@4dor(�1!Z�Qwr���rpIʃ&���А�mM~8R�PNֱ Q�W�&��e�̀P�$.�Z1���� 2)^��%��&�ɑٿ��þ�)�9̠�3t�.s:3ߠ�L����#���L����`n��,j�(���jD�N=o��i��&��������u��?ÇfE^����|�+���e����7f���Ьm��aV.,ڒz�	I����!8�G�%P�/K��.���ǧ�f��X@3H�×?O$ן
��g�N��V^��):�`��k�1Cn��Q�!�[�Ie1����Z�=��C��7-W2��w;�-�6?[��0b߮Z-�ƄbI����|.I�������*q���=S��w�d�_ћ��>���>�Va�OJ��ă��k�]�zJOЮ$�<�U���H�P���L����S��P����<���9x���
��`�^4�z·��9�,�DT��ekq�%��a�!��������*�b���My	�S������;��[C���b�g������jH���/��c�8ėI�&���Ya���[7]�5J@�։�0ݼ|�Y��}��S��t?֌���*^��%��D����p+�s�1~�1��� �6�	��OV�'����G�Sh��s��B"�J�Z���,_a�[�~A|RMC��d�w;�!�.Ԩ�`E��Ӗɣ���o��B����\tĄ��:�m�!�f���#�@V���,n\۰tFx�Ⱥ��S��q��=�4�ۚ���Î�,r�6�v�mu]����Q�e:���~�܋����0�>��ϣoW��`&�ڛ�Y��/n�X���&���s�xP�w����(���,,)PG�+b���#����_"{������aP"y*|�Pd#3��U��YUo=yu�t~|�(�O�o�áq.x�N�A��y)����ה�;�� ���IA:��󅋿�^��]�
C�ߥ$�f�*ƻ,a:wɖI���D0n�����7�07�Uo|c�#<��j�n���;��m����Xj �s`��tJ#�@���տ�M5@���$���,��Poֈ����D�"E��Q�x����Mk~�DЋ�=����4�Fx�S\_sc][8Q��$��" =�"Sg�٢Ll�I�ι��ǎJJ�ٷpFc��q+�5�Ps�ED&`�WI󡿷5ӄ�b�y`�����[ �<@Ġ)�\#N'�2�nyT�*�ӭ~J�ۋ��aF=�{Rx��|��r=�U0�Q®���C�'uN���ޞ��a��s]?����>q���O�^�x��P4��������eK��F���o���ۦ���k(	L[����9�;L�RMg(�v{}��Q��9���,~)�j|�ksA�a�*��!��Jp��Gyy/k��ڹ�ٚY�S�8���.���Gf%�dl`�s]��g�V1<�j⡤�<W��u Ŗ��8��lbE�����74~�,b��?}�A'���@�F8Q�Mv��Tq��N� Ce��N�#-��[J�>@kgm�Ҹ��z���6�W��TH�Y���ɳũ��ށ�e]Q��c^����ip�}uz��a~'Q A`Ho��3:�A��e��G�w]i��>�#*�IlڏRR{ƇOXk [����-;,͈o���� ��3��,�\'r�����8�)1����I��|����힫/�܈�,G�*J���k$s�h����"�n��V�wSzX�)�T�����v��\������B zCQ�26�tJ�-K��O�r�:b���s-q�W���S��x;P9Y�p	��`i�a4C��u_�;��-5�v@$Gd:�U脤x�� {2���g��.�/et�G�]�T�ې�ͪ�ih�-|O܅Ar�Т��!����\dj+w�oqɶ�ͧ� 2���pm��$f�.l��o�1�=�80m�����|
J�
�GN�� ���7/��EM+L��^h��_��>��Y(��R�)��cbgԻ���}>�m|�����=�'��`��m��xE�I�F_ͳ���˱FP�=Ԙ�2 �s_v��#<ԛ~�^h4�o��T�V�*�?�Iq�!W�;'�Q$��ڐT�5�b/,t{�n,B�	=ۺ���e$̎q>���Ѱ���G����|��Y������Z���ǣ�w��w��i��h�ȴ}��BIS-9�{��y�B@��L�R�x��7�r�:��|U�d5XlxVHYEB    fa00    1d20kFF9*�a(M���� ki.ʹ�=�TB�m-V +M��{"f|�bR����!x�1S�Qe�a�$�l�8��3	��xD��u��Ǖ���G�[a�Ȏ��H�mт}i�T/��I������������x�o8ԅ߫�0߿g�Y=���#-�a�=G5��($L�f=�2xT�9S�j�Q��d5;� ��M�}Ou#nw�B~�Vw�r<2s��L��F���U�Ȣs�%9M�n�S�^>�r����Q(����yɞ��oEλ�]ʛ�/����p�2A�6�~:������>����n+k����F�e�j#�ŉUA�B������D�ܱW�&�ؿIg���kۑ��|^���L�gM�bv�t)��@�gނ^M��[���k�57�����yu)�_�2�M���vGq��=�x|��ˏ)�|{��p�@}xn���&�p�����S�>�znn��l���EZOI�b�r[��t�"<2��T~���( ��B)��+˩�j��[����n_��[�~��Rώ7E��/ 2}�:�?:�ۚ���+����^�{t�ћ���+��To�z���T����ˇ��.��bt�R���6bB����<�6����X�8)C=7Zz��;Qn��K�(�*�i���5$`�� �����w�Y��[O-q���J�`��
�f?$�(��U�/�?���'V�;T��KEO�˓�G4�+���{3�ra��5�����s,���Z�.�E1����x�y��@�-,�T?+=�a!l��6�gs�<Y��V6a_�O�Ik����4�t�8���J4N��d���G�'�'�X�%KxE�-]$����â�>n�I�Ąշo�D���.o��L&�پ�@d�ffX�3�]�xG�T���t4 ��A�u��O"����o��|���KǠo3�k��z[�ʚMZ��.�f��b�mwa�iV���	k*�VH"κ�#�f��N@ 0�3Q'��]ۓK���N��Y���r#_�a���eV�j�.� �J�[�d��k����ӈ^���W����p�/�Z�ѯMIf�K�{�^�d�����ђ_4oY�3d����J�+h��k9��W��t��2���m9�oӊ$�Ww��B��/](�4R /�x��8�ʑUތ��
�i���Kz����Iн<��lR���eĸ�0g����+x�p\�����l�eԮT)���vbζ<���W-��I��4o+��jmCY=�U*>�W�~��w��i x�z@;���$#e�!&A����00]F�L��)�Kb�;�Ҩ9Zo�	2ڞ�4��fk[%�Үn�i��TE��ۍ�H�b:S�<R9�\З���2�c˟����/���Z��u�X��p�R���
t(�ۜۓ��Wu�P���6�:�Bj�����0���?���Q��=U<�36$�5L�%��}
�"���/bMY��o��4�.�`���&�N�?�<R�r��C �S�r��x5�%�B��~ظ.4r�
=�J��/$�P3��|�m����Z���{����R�Ak����+k2��KH�#���h�t��d,�!�ր�}�A�l�=�����M��a/W���	| i��*ڶ�/�Ts�q�S�߻�hu�mJ=�P;�:��>�1oBAB~>zڄw�0�4��$e?3%��ڤ%ҳ�}b�+� =$y�H������s���j шV�������ᾉ�br��$���t*�����7��I�gܦxဇ�݉�c����/��Y����p�R�.���f�ܣ�ٚpm���h����ۀ�%�#�}D3Kl��~��_��� ����s�Yi�mQ,��,S�5 �
d9���HA�i׃�H�3��,�d6�M�ꮲV�ܼ���20�\��B�5P���ҡ3zH��2��n��ù�ܹYf���.�9ɫ�~)��W���'|��&B
�CY�Q�uE5���������X�{=���k˞�eԨ�C�n�e w�O��nI?�JD1�I�(8Y�kT�P/Ս�ן�l�І'��%_.S?M��i�6�^{'a� WJ���$���9~c�$ȱN/v�&�ɽ0�1ơa $&C�2�N4���4�����t�fcc0�U+#' Ȕ�p0�#��*�^P�M̝�,�N�N,��Τ}����X&�O���|��5�$nPB�/��:�XEn(�����ǎ &t���"�<e.��&D���tO����2�祺Ɂ�4ʰ��iH��Wt�"V�r��ka��M���%�~�,�R��i@,����L��^�7��M!�R�:O�������N��.�=�Y�*OҺ}4}��R��G]��К ���F֟_*P]�
�DQ�8:��ޝS$���T�O�=X*m����Fy0�
����\��.����(@	I`��˹bq��f��ıТMh;�W�C�X�t+:�%�g<���2�������|-�2�Vō.K9K'�: �l7E�/ئ�NW�}s�2�"6�~��T��躟�F�����vz�RPT9ƶ��ݴ����#�и���k�(���"gs/s�mk�(�_�]ߎ�:�,^�&='����Q$a�L�I���KMi�eu�5�4�͠�j��� �,"�j�j
iJq"o����B��_��k���ǂ"|[�@άM3��`E�1���M����f[^K�8`9�P��S�f���̹��=��'|��ۇ�=B����$Б��KE��zm�eq���=��)�kЈ�\I�c�)a�EQ8B����($�LP��K��E�*�۱�x	D 0[zs^Nbw�!�&�g��;�vw���V�ɧ}~�I�����Ԙ��O���u��/TB�_On���1�-�ƛ�(r�z~�(A,�7��h��P뱊�pȊ�޽Y���+�x�ud�}��;5^�B����[��~����P �Ύ���Q�N�}���ث�I�ddXX������F��l)�R9ʩ����tI��n�0���I��"P�K�u��340Ⱦt�ǶܣBri��)����7C���@�4���MP�bLu�1l��%B*�j�=P'J:�gpLa���&PM�v����$�mi��R�IN'�p�F���/��>�����;�������^�qc.�N���5C�|�\*���7�4\�ًo�g���׽�(OM���_ެ7�&�|��0�]��)�㒂B1𬚨|P�B���%����a$1����I5{L�|�������i���򪎫��Kc~����IU�'�R\������O�@��ϓ�{��%\t<�����cG�(��[ӻ�h �u������&�k)�"����=s��rZ��#a��|ǜ�9���0�dI�����]L�⇴<�4w~ �6eOn�X�q�i�T�%»�E�Qa(���*b������?j�bN��E7O�g��$(���a�>��R�40,uɷ�6��-��l�"�����ץ����q�g�d�h�*�w�J�����9�v�N�?�%P���E�	r����ԛ���/����C���l���gm�eQ��>��@Z���'!���V^=T�rZK��8�Y����A�����X+`�<_7���:,��#QYo}�f?�D7HSQ:!ў�X�-�a�9䓨��۬]����Gb������@�j*���n/�	�À��{I� _��ǿ��q0W#O%Dp��$�I��l�`R�md�C���,*Rݍ�l6�\���7���t��0V�Nd�ы�{��v@���x��D�ծW(⩽=0&��q���E��1'ߠy ��|(���>�����mo�5;7I��AAJ�}c�!GY���MB�E2\"5��O_�1�>�s�uM��B" &a{K>,X�Z�x�D�bb��y�C� �s�V��'��劣q�?0��}���r�����9d���|�{�F9㏓�E�}�
�F�pt~[�ȩ�[�O�r,E"X���-�ū�X҃_�3��cYW����Wb����@Ϸ�BzĢ-�>0Ny�J�4���`�����޼��J�M5@_�MI�'���T�6��õ��ȃw��N=`�|ǌ��˖�R�Z�E��u���\±w�&�m��%w��j��!�l��*�c��ub�n�$Ͷ}y2q�����_�L'�Bo��K��O�@�&I���ƏQpMa8SQ�������~�9Ҷ;b��Q;/"�0xjn�I�������fG>��m�⤜��`�V̿���
��%z��Iw�	Ӣ��ҒL$&�]� x���}��΂�D�b�����M����T�bؿ�Qu�'#4�l��t���/�mZ@$<�g�>n1*�Ȣh�V|��n�i\S�X�(��З�jxif$J<��h@��Z��5��j�]�<iOK� )B� �8q�n�ܶ�����ѹ�Q�((J��x����"͞q���ܭ��C&m���M;i�Z��:MK����9�'-��g(�`��n��L[�)�9�.݀B�U�`�1�$�O�t��Lf��'�|p��݇bW��3c������;B7'V�n]���p�ˢ��1:y3�0K֋�ܑ�yL>�Wi��	*�1����@��v���Ire5Q0J�:S�[��-E��%uE�f=���>UT�"T�>�twT?���`��f�C����Q���i�ͭ��nMӓ�~���%ܤ+t�hb�=n�	p%�u�>���?���27�ɠ<x<���R��59A�(��ݵD�����.�(���բ��.���n�K���*�ͭ���jt�[8�z��?B�c�_}P�������+ωWDf[�7�]��&����(�����G���h�V��o�i~�hϖ?u�"\��m�Z,RE��D�Y�\�eb���M��{12
��C�_��)ۆ3�U��~G>@]r()O��"�^���ODhf�E_B�x.E÷�T��Nm8h&���l��h1�gö�_l��ܩ������{�U���/{�	s�|�O��%�N���y2����Uv�!�t���?΁�!6�¾���,X�~��X!�d�jpB��X]�B{���ѡ�<|^�c��H�����r��(�f#I¼m`;�2��tI�!�6fKj\��]�����ѝ�Г����@�������B6 T�?�O:t��'�����3<�1���&����ke�,z����<FbN�X '&U���7�E��J_���\NǖH	�Լ�/����ƓE%�S�ұ<@��I]�&�^ՓB�&#3����]xI�F4����e����R��KK�Չpx�ǆ�?񐊯��7"2�\=ơ�K�r���@����B_�}��7\%�C~�jo̷TE��s���2׆�G��3d0zn�2�+XBu!�np	��*����(᳹U��̡j��*0|!� ڜ�?���9��YqcC�B?���?��� ��@n`����e�o�K�P�;��A�A�(a�LV7��e�J�R��gNU>m�~>�J��M��M�H)��v�<�C��<�����\��Ӓ�L�����QU3����"K*mU�T�,Q�L ��� b����0	���-W��>ٙDf��SA�/oaW=��=L���{:����/x��������K�DTT��� V��$��`)̎o��%�e�}��<n�.��Y+@�%�`.��njD� �*s��������h��$I`���晤cr��>'LN��q5'Y��a9A���������U�c� �j���Q�|[{ٶ����鿒�R�$ۢD�l�N������][�W>����?��"_�Ղ��F��7����՜�׈�Wf���t"���8�(�����'�t9
k$�;��`kC̓%�$�۷6|7�I���Ě 1�d1��r�������)n�n �Y�E=9�pVL����(�
<$��c�����I'�R�7�v�N��'=���[��}���;@�È����N��@���݉t7$`�W��?���:J�	�B:P�����y�[���(*���`�>^����� �i��ǐ�!���E���dBn�1x/�J�����(dQ���;+ss���g+GQ�����w'��1A�f�K�:��1M�}�,�~��8����wA'=�0�sq�;�h�	�F�(\��ŚdRs=aF��/�Mr��@�%˹Y}���>��J��9'�얾n�N��%����d��_�NS�i�l�,{��]8etťwˮ�G�KX��lB���E����H��7wN������D����'�|��:�χW7B�����"�k�^��`�۵E2��̽ �w�*�xk�m��\�/�	��f��;Ҵ?�GyxXn���câ���d�[ա��H�6��2|�\�o	1C�US�Hhm� ���H��W|�)n���2Ob�b�r�|2��t)qF��O��b3�#f���E\�ֳ\Vq^zHrC�G��N�j������f����w!q2M���{��'�P�N#���r8B����G����ҋL���6=�h_�g@����r�`֨xh�j�#��1��'�s��
T�����S6�=0�Hx],�e=|
`�W\(���*��Ja����z%c�gচ$�=0XD7ڤ�_�v�Y2.ރn�[&�-�kqG�r�;Yݚ�Ğ~�n���]��Z�LD��0�d'6:h�ᥣ�����{�`s+�� 6t��x�4�#Kt"{/��Qy�3S��K�?���@ɤ���u� ��]&10P qY6G������,�-����鷤D=8i�q�S�Me�%�?��m��IZ���\qn��L��n3MO�����5�G�d*LG�:��}9�X�G�@z&�M�M� �WO��m�y��~��om�'E �z�Y��b��Z�Y���/�Q�S
���s�n(-���`HB�^��^�����y)F��=�d���W�#�(��(�h�n���s5m�6����b��%�Ĭ��(�l��s���l}�ě�fa�C�y����l|��\˲\l8e�ՉTjB��(��!s�y-��^j�S�d�։,N�T�Zk�[����~���t�=��d���������e�|�YE!�k�Q�۹P��1���`�~��/J�@p������;��Ǭ��t��h���R�<?����3�́~d�I�\���["�О��5r.�g��i
;{����B0SΤ{���^�iOZ 4��[(/"9�(�����G����\��$UzPy����m��Z�>��vn���zO����<��"	�����w��E"=)��h��iF���PP��Ȥ�0XlxVHYEB    fa00    1e20հ:S���N�Ҋ�N{�G��Y{�Ċ�#XI��29������"���>�#��t�y61\��Xj&",��OO�NR�֮�1."y���Tr(HO��@M�ݙ���)�C�ǎ�j�&v�����K��o��7єo~�!pF=��\�N,�U���NE�
�� ��t�vO��ʻ�oV��p�~L��E�)�_�l�&� ���n1D����T�Z.�Oq�X%����ߑ+`c��s$جy��k������h�o����E*��3���4D����<`{��
am�� ax�x&,J�n�s���tm>�ht�*^m��}�C�Y���E(V��.U���d�z'vl�
�����x����$t���a&�q$BkԴ-�����w��2_�$���3�Pi#�971��zBcC&[��ůE�wp�B�~ܹ���=����U�
�ߨ�04��c��AɁ^�-ۜ�:6Jv^��{�[�K�c8�#!R
H�e+T%���@� KC�����bV�Djz��E�҇XR��Q��azѯb��ٴe�\�����c��6��Jq� ̝�b�᙭n���[�9�U��]���Cы,�dm����\, L�R5�)�4����u��(����ƻ
ߝ��i�aP�+RV�1EQf�F�YQ��^b�d@��H�|Xb�(��/�.���_4����R�t\t��w5p�[EZsn!��d)��"�q��rC��F��-Ǿ�$wF]���Wst��"�3n�<�*43�[jDǹ6z�C�(|���@5#A�f��Z<�h�2����D*��x'��S���0Cn�M��:L@pӜ���^o�[�sSI\�7{�]�D]�Ŝ�E�bs���oBd�F�)-�(NVȩq���'u��N�U~~�*��NQ�{��� �.�I<N�`@�t�����
ự��`0����%3��]�o�/U��oi40_ ����~L�f��9
PC̱=ܣ��!�������2q���s%�#f
˝�d�Ũ��Z���D��8��J�9ly�'ÂJ�4Y��$���ļ"�I� 
��k�p��s:~*H�n6*Z<�لE� k���ؾ�-���-?2��Ҵ�]D����V�BX0~�0�
2vНF+,~F�$�ԴP��D̀?�$eA�u��>1��s�H9����7|�6+�޳�n����& ~׳쩤�1�@\�N
��^ N�tȸ7�N[�%DM�J	V6w���t�H"��1g�d�B�'�SWH�DQ�������|"��R\���N{ô�/�/n��)d{�"�#C�Sɔǰ��So��2&'�)�R�y����5��i���U&[lJ[=T��v��$5��{qF��.�G\�q8�yH���FT�	vpr�ҳ�7�,H�b��}�&�쬔�k5J�B����v^�EX�<�Ry�	�7��`y��pX?<���#��6���9=|@�S��J_����=쮆Ͷ�Seu��\x􋧛x�g�ɴ-S�:�^��CFʻ�?�����f`�bkƋ^�b!9xrV����Gm�<��6�A���/)�H�����Mk�a���i��eЉA7�N�|l�}1�H���_���n��',Xh[n��K얱��>_N�ki�ՁjB��Un]���D��K-��^j�3ʓS�N�����N:n���I�4K�;7�0��Be����I�T�0�4^�S���l|#���Y��H[�Eb͆�6�n�����v)�'Wwg�U�?L
зڌ6��f�@J����J>*��j���~���f����).}?����*��X1��+IܕJ5Kftkb�a���D����aJ������l!�w�`���Ũ�u�=ϩ�G��Uu�dc׼�K�Em/|U>�Z���)��x�f�ͽH�C���+�����~��^�m��Ri5��������ZdX��4�#�[;�� ���d!��x$_�7K������� F|�A�Y��0u��;p��i�mr�3 �� y��HG�����fl�� y�gB�y��_]o��Cȥ��Pf�&}�k��_�* �-2�{8��4]�<=̡�2;�
�x�����d�GX������G��y�M=�oj�J$ݷ�xGU=�@��X�C��%0|���0�:�E9f5̈́;��e�3C릺E��Y%�0��l ���5���b��c�4�kRZ���/d_��x�	}��xq�*4�I��<�ࡉ�A�E���TDm��g����vCL,�5��h�r��C]5g�Ʃ�6���QF*�zHph%̐�j~�1pߔ�a����?�L56���D��F��:27�l��/�&�e�eC�O�/���;c����
����/�Q�%�9���s��.� H_G���'����z����@3�����X{���p;ꤕ �I�3�6�� �k����\��*>�9[�pO2�b�E�նs>\�t1h�Ҙo�L-\\j諞�sq!V�c3�yr����X0���g���@�}����Lg.��Rx�83V��rK[㬎�iS������>�e��Q2�!�_���&pJ�,��-���f4ݢ��ya[���S�i�%G��+jv�ZL��TQ�,� �Jv�, ���k���e��(���+$����|�p�̸t�a�@�W��l�t+�]���ƪq�S��A[賈^pQ������%p��5��{��7�G$�L�W��^M�Pdf�C�0X��?qB���%����w�S�
���R�v�+T1W|����B����gS1&�y�� ���.�w���?���ޑ����z^O��ot&ʰ4�#.�<%̑4��s�� ѳRU�7����ifuV!�T7�Z�`8 Ho{�OH�,Ug��'��}�N*�S�j��W."&!�x4�o�V�Z�B|�(��)��7� Q�+��05��6g�xg1[��nzU�|����jW���v�@��18yݪ��n7^�5��W��ٜ�Ƴ���ss��/�N[������Og��;�S#�u?,��B�~�ߑ��Y��B�t&�`��:<�"*A���n�Y�n�VL��n���f���`�j�����qJK���Y� ޤ Z�=�=��tW�52�C�
j\����t���ђ�>O�V�Z��~{e��f~T$��dt_���8[�^�_�J5m63�nʧ��W�*IlS�*oX��=�P���lYmx�@2�H����OL.�����NWx�zb�p�b���iw�^�Ꮴ��O
^d�{�r6����P�q����i��n`ԫ��g��������[�L�J�a�%R7O��]c�}�u]P��$�ɕݓ�[�;`�9���`H�y4��q�9���y+��/��3�-����� #����A���5gv�4~H�A�8n-!! ��S���*� ��lo�4�U-�0�Պ�q�y^�f�`�XW��	.�;w���ME$�$�z��k�Y�Jh��}��t����O;N��� �}8e��A�@���?%���3s�W����Bgĝ]�~6B�g���ꙇ�����i�dc�Iw�!Ֆ�����wK�q��^�dg�F�ߴ@8����*_���Ys��(��Q�\}�^��-]sD��l#��]��_�k,(zy�>����E���n���#�S��Q�I:"p�'
��4�l���?K�D|h>�;�yuG�&��%����OY��T8�oi2�(]`|��E�lu<|;���g5[m�.�U��&�*Ӂ��� M{�XBm�LոB��_Eu[�&;U!�X������Ni�M�ٲ`�7$2�O�I6E���!�ҋ�7+�vVn���b�'i�<����n�J�����]�c�9�X�n�(��4	���1��i��dZճ�����RF���w��Ӕ���3X��·��B��)*����V��*�� d�UO��"���aR�D|.�����8�������P�nR�&2OҨ[a���f����د��A�u˞%'��-�6��R?a�(��E��B=)����@[�oH+ڄ������N�
�_,,ϼO��]���uKzY�u
3��p�?Cכ��Ѥi﨧{�b��4ދ�hf�FA
�_M��Վ� �0��N
��������+b���YUɔ���=ZF�y���i��%(�q�rXu�e��&�h#To��>1`�}S�\�8=�����3����8�@&�.
OP�JU�u�o��7�`	�n����g��^�j29���&������֎��i6���`��@�G;����,���u��0�n,$��K���Bt ���я�w���8�ug3a��m���|�nilS/b��hM��e��馸X2�?�"i?�������zX@����[�+���x�[�z�7��?RT�2s���nGm���A��iV���ɼ����^�M��s�A��h�ej(��?�z�N�I4]�`���^�F�8���:��?*�y�n+>3M;�(6$��,:�#˟ �Z��5jd>h@�Sرm�͊�P#���\�z49�.מ�7({E�{����3�b���v!n�JPG/����֟��)�����h�-����D�8�Iz⠲�⣡�Ÿ�I:�����qr3Mh'�=�o����4ש�O�F�U��l6��2xOG�0A׍��<ۼ�BW6j[ڟ���~�<�{�ꒀ�rR������&Rq����!.���t�O9O�2x��Y�|�'c�����͊�J��;<��=��.J�+�� �ꀸ91,��9�؇ń��v%�<�.��������+)��=�[}V��mHW���ly�@n!�&�H�$k�Y���9ӷH|�\7M
�!�; @�yN����4Hw�j�?+<c�A<� ��7�������?�P��iw>���M1�Ib���%���[tG	w^m�a�(\�z�H��뽿N��!�Wx�1 ��q4�N�ä��o�BW���`d)��1������[�L`�21r ~a+�/�2[Y��������N�&����~���M��)�T:�$��TƢa����$��G���	�-dI8��n���X7�PF�Is�t���{eg��nw���-��2W��.nfAjکt�n�A>3'&�S��n����m������0�����ik-�{h���[_��M�ϖ��+�3[*��z�D��9�!�lS'�K�v��( w���+e��<o}�\C�@��b��x.����0��;sM�/��rgpyE�ST1��o�]�� �/���ϔ=�b��)��q��+]����^�t��׈9�y��h�%j/�!q���*uW�Ŝ����|�A�S�HTH,���h�1�\ �� {�����_���o+�EYT��[C��P|R�'�F���0�O�9i�Z�=���آ��O���)���A�R�R���>V�ֳ�(���N��}�	���Mm�:��c���=g�c��M���ڈ~��������@mV	6�دޜ�&��-��$<Gʗ���0w|x�G�!P�퉨��HV�M�ohAj4k��t�pUyB%�,ڄ�I�"�
$�,˲y�K,��Hm�If�Ry�ȝF�m9�PCC��kR5��n�k� �ڥѕAu3U����$u�x�&*��R66���M��Mmvښ�j���&��{�sӰ�xX�a�G��r� �s�~Տ�y-�)�T�e?}�!�V����T�T�>l��r�Nv���K~�c��r�{y7t��F�V9�b+�S�Uy�̧_�r���T�gQuU��zZ�Z!�"KП��5�������a����i;!��s���a����fݡ�͉nK��D[����7�O�|I�����_�8Z�4��wk��̚��}O��0���Hp@�NsH4�hX��9�q�F�V����	��IO^q]�}�5���߆fm�N;)?N�a���sЏ����DP�]b���y������s*�$qa�2��$�8a�&�Ψ8�z'�4�Ur
�'iA�@	۩c�ȢV2i���ÚK-[�;il�[��ڈ���(RJ6��l�D_a\m�����|MZ�uRg�����2�����r���8��WJ[�7�*��:��,�YS�0LvM�� �xޜ�l�|��}$����s��mٗ�BOfB�W+���Q�c{�;)�U�#9�"v]��x���#����5F����Z����?���]�����j��+N��^���ɹG#7y{�����M�02E6�A&�&f�\t$妈˰��\�;P�G�D�}����!�ܳ힣��W��)�ܧ���,ڻڑ#i�YΊ���Q�C�ڕ�������vA� P�K��	q[D-�;r&R�����6��#T�ɒ���s2�=�P���� uZ������"�;�(⡒�>O���Ҙ��l>d'�.V��:�rq��T���1^5��@��"U���&���+�%�7J�6amiЀ������m�;>d�W��l勁���W���گ�Z#�G�m�8�wݰ�> �Z��ě?L�%��=�*��B�1��g�{^Z凮s�u7qE�:�:���x�����g��ڃ�ߡ�@d�n�s�F��� _��DW�/�L�k�(����-Į�m� �f�������������r����xK��/��w:�d��U˒$�
�Wr��x��w,�����+���;:�����a>��"��洐e��-@�ў���b�4�o���'���N� �8����L��Q�v������,[c�����a�N:��Dl�ڱ̨�ggq1^��j�H����%z����d�7N	����)u
a���)!�v^ )u�}��
3�0���c�bK��O��`uOG�$�T���3�O�~�M^�H2��b�� 2�v�&EcM.�x�Pt�w����&��*ob��}��(�afjR���_�K�k�;u���6L����OSN8��ke
��V ���o�WB�TD��	;P<�+;�F6C2nB|��t����F �+H�Y�S��)�>?�a`�r�k��ƒ��=����u�@d�ǯm��4��"�v����J��'�μ�8�ocYCz6T�CK�y��l3�8D��,�4p�ɹ�'���)�C)pݑ�+LL��\���GA_qȹ2UP~�f�&3+p�����T����|�:$@�����2�%��xO��)���LE	DϞ3�mp���@}&������s��Hʤ�&���˹���J�448�J��Ba�"�w��Z�`���0��_CaU��ϪE6E�4+���� ����F~��@��ho,;�֝�|k �uI�Qw�#�r`6�*�Q�W��m���<�y��%H���ל��u,X��~R�j

���Ԧ^t��mn:6^�܄y�U�]�i��3��6	��������Ze|F�Q���P�;�It������N
�q����½$�ӕ�	x����@I�/����1Rx�3��cv+��r��=ͤ�J2,a4��k��V����z.=�0O�
L�#��+��	��U��;�J�1$���ǎ���m0���tv�5ߜj}+�e�.�bX:Ɍ�)S�ֽо=�%P�D�� IՂ�2.F�$���W?�ʝ�-�4@׉�iXlxVHYEB    fa00    1e50���T��X��3�P-��I�����޽�pb���פH�A�O==�����̴J���Lq�����"�0c*M!H�%�7�-��R���e���PvV4$|�TE���Zڼ��3����ߤ�C�'���D揬~���� ��^E��]��QI� ӓ�����!C�L�R�"�LEЛR9D�L*���B���Seţ���5�r>��F{�HnX
7�`�Rh������l�e�+�>�%�-~� �h3��Ql�kO����&�@}�bb?�����6�m��Z<c,_Z�=∾���ٍ`VU%�JMf�bc%z	���A��  �D	2��o4�/Sm�5qd�
D�M[f���gZ�L��H��$����W7q,�B�M�N0q�x"���&q��4j��C�a��9q#*E9����W�RM[e4Co���=7ci/u�I3rΠ���!��u�̺q{o'$�˄���?9�*ۭ��2�;����hJwE�<䨍J\���8M����V0c���R��Sk9�ө��E�eK��w���*��/DˑnN,���i���7
�T!|R7Ѵ�z��D⤶ŷt��|v{��:8�r��FSy�çl�m�vb��i�!qj��q¢ez	5� �pr�D;�YW��oo�`�KԺ��ɅZ�MC%Y�K!�����{7���`]��i �n�:�[�«�4	\��Gj�?`|�O4�H�:@����#���γ|&��ʣRZ8��JĜ'uG���aOUb¯�C�{���銾��ð��Py�p�x"W�2��'����J0�C���,ڞ��gtָ28k �&Cw���O����M1���e��:$�#��s�օa>�
���#���-E��hvJQ������8?�U%Q���H�O�`���j���wsJB�o���e�˕	9�W��'�&j��|�6oq�~�Z�l\mABn诱H`B��Ӏ��-yu��;T� ���^�)l?����n�wL"C|���ţ�Ej�)��&�ٸ(X8�X��Յ�%�x�A��a��2�On�j<M�/\�]�UZ�_��������TSS^��X�^�QTzh�B��� tR3�a����_���1���2j�V�Z�w�(vJ9*j/��]�ʂ�v��ە�M��%�Y|q�r|[U[�^�Er�ܡ滷$+�$�p7�E�cPڊ�:�����\�/.�c�������K��G�ęK�y.�����O���Lҏ�:���p�5�5�/f	=���;�i�0@=�����'=Z�_L`�X�7<j��Gɱ}��ی�E�P ����ig)�q���ĎG�ŸEGHO�ح8�gl���A�g
A��;&|u�A�H��W�}�ov��}�0�Un��QU,�!,V�n��(_����3+�]3�x�٪�/������G��j0xp�$ƥ���d8a,��D��UNAX��[R����7��t�٭ Ws�pV^轫�L �\��gŨi��?D��B��%���$����C�ӜE߲��Wi�aCkan^#Z�-��Y�a��12�����w�j�&mn9�CyD�^���&Q��x���C�*3+��nK3�*KX�z	œz�qŰ$|��a:���%�N[�r	.�
6K%8����i��{ �Q�D
�?�����pdЬr�=us�i�+t��``��f�S��?�H��
	)$]���P��AtF���ds
���_P맅�fq��\%��t���u�!:��3W��?�U!�N����2�s�j�xa�К�a,q��_��t�Ȏ���*������1U��Д�y^%n�����?���|I�}j��ڗ�Z��N�UKd��[3Xx�i��p\՟6�~��PO/�&Gej�����p�}�y.=�-�9��V���X<�0T`�X�)��G� |���g7��r�k�Ɂ���L��7ե"N�_N�P�k,K��zö\j��gx�W$���!�.�W�!Q��zN�ѐ#�|�$jIr��=St͜%}o�!����4��[᲻�wa������c�][�Z��j�Z�e��.���[� =o��V�/����G|���z)$�In�z8_qT��] {��$�n��#To�(+�?��|�����"�� Os�h�!tVs��j��I��%����[RT�u�o'��K���(&)�<.o'�/ǹ-mX
�+Lօ��	[���͵�����`A�b���/Y-+�7�Hf����C�/_���)"���Z��m'�湯�,B�[S~�m��V�`�pm��7E0��;J&��Y�I�3>U���u��M2&^�3$���ژ̰� *z��q�l̚�Oߞ���Y]sN�N��:����ٓ%��Z<�5  C�򨤝��M�������c����#~��N<��1?�3�(}8�Ogd��3�43,R�-�k5��&��CԚ�Ͱ/"�UqRz�`��F=�B�^�LN�TxP�P�H ,��h{���J�]�2�6��)�ˡf;)#��f"%���
����,+��٭����r�������J9:#��_3p!5������:��Wh���6����u��!�֜����0	C^�־�_Lk�]>z�տ!���BbM�ԋv�*^���_u~������0:�{�e��g4GU����r�2�rWNI�ro����~���@��ATP����Y~C(v-6(�1GP�|��rt�-�|2��If���� �6�E9"���$�P4��Tq{�D���L����r�;�i�zW�����!z&y�.����w��[�6g_����$�C땥��b!�M����*�RaW����y�s�6	� )|��ɹ1����&9e��/N�(��+��U~[��k�a�R늛����>s��ͬiE;j��p�z���"��҉DDd����Z�*ѫ���N���u�0����E57=�o1��P0D�61��Y�ҫ��Yk���%"����s/"2�i�G���C����R��:b��@�J���6���|L��ŗ/)��	�����Ƴ��u!U�"��X�CǺJ����ު^��-:�b(�n�jp���pW�i�Jq�	<��PڂⰨ��Y�T�K��V�f"�^/�BF�)�n�U��0w2���d����Y�c6�lҁ�����p�ə���V��0-\'�Y�;�� :��'�#��Y%��	f}|�Lp=/�r�PJ��pq��2E@9���o^�8���t�Y}c҉qI�Tu�{Z8���vB����i�~�D<�-n��.�,岵�dE>ݙ&���Y�39��Zr9��Y�1��;�q�mz!��X��و�.���b�V��V�Y�.��\^m��|�ʑ\���=<��5�����%��ᥭs�j���GG$��8������Op@�sqK��?i�{A��\5�K	����@s�Y2���u5\��^h��'rm���'����Z�?W��Ϸ�k_{ǻ@���"����k�7j�lX�t��Gs�$��	)8' �Ql���[|�c��$����;F�@���h��*!�UB{r�!@6���W4�s�'*j*{�Ù
��i��F��L���yda�
�{.�ɚ����d��9wSV�����]=����Z��m'T� ��)We�Zl�'��%n�%�G>���׏�Ӡλ;|V��a����x\����{��v	)�F�=�wc�Hk�93Ħ'ř@i9��GD����Z�ޘ9��ye���Nn�=����\E�Q��r:����4��h�[\��4�{���cՉ2}N�'ޓ֥&`������3�H��k#�'��1��6	��;�0bi�14�:���g��T<ɓ>P�m#��H���_�O+ۅ����^U2���r�C*K1bN-���0|��AJװ<~���M����U� H%�V�HD-I=j'C��`�b��LZ�J[��\�Iu9��T>�[j�e��<=M��cS�����qg-j�17�ק
+��f��*�lc��?�Q�B<_�����t:�@e����^+��Ճ$�}�O��,�3�DN:K`P6"^�-��>�:��������&՚6�	f9O[lp����G���KS����ӼEwM%���ux��
����Em7Ȩ�#�}F���:�T�EÇQ�U#������d;�b��[�ñC��ֳ��P��׃�8�cp�G�r�~s�[�U����4�ݞU�D5ʨD�[8��t��L��t�( +�)ǨM~��+�~�����.� ��&�佴X�"qU^R��q=<-[�;��B��I��ix��R�$f�ݞ��y軚��lg�ԏP�3��9�."�#h���*�vn�\�`�ߜ�*�/�l2>�ݽ��y�ж���q 
��jω��ǿx��T���>��
�\Ր��׀��<˨h :��U�`OOC�>�k���(���s�s�棣Y�f<�'/�I�Dz��4ս�,)�KdD�?�҃}T��&�ϥD�2�gv�jý	���6r�Va� 502���ds���}��JBkLo9+�P/Bo���{���k��Tf�Yx��%�.B�/
����θ�{��x[��әdµOm�:�E�q�`x�
�v@U	B�iU�!S]��t�i��(�%$�?t��Pj�4�DrAݛ��%F�F���W����9�ʟ[
D���H�b����d�G��6���p���-歰x푀��x�?m5�V5��W��,�p��O�c�I��]���!1��Dvbś������h�B�,f�kg"F���Ǣ�+0�P$��,�K;o����a�6d&j"��|��XJ��Ͽ����c���F�b*;GNd�}�:z��G�sb0FD�ei�O��Ш:��=���5&^�[�KU��t�C6;*��Q mJ��X����R,6��W�`Be��L���Fvq<�s�ڦ�$��j.kN]�9�>�:{��_����p����\&pf�d����t�-�Чcc��冩Y�r�D�5v���j�!C�&ya]T�V��_�:�K��^�y��;�{�~KVa�O�?~׾9�=���R��3E�>ܙ�Sp�����4�,Rz���|aj:�w_@Ӛ��]ԣ�s�}�5�ug'D|�;�f�t"��@�6���WʂG�p�Ұ�t%�聟��Sz��Ujf��ɨ�Y�˗[��1OF�2*u.׭J*����E��]�)Ɖa��G�Wl���`��2&�3���A�gXT|���U@۲����`�?�:��
�
o#۠K���M��˄S��������ß��<�>v�徨IQ$�SIix��+�����W2��M(�lp�+KFI.�U�F���$�1���6���$+���J������l�l&יŢ�>qO�'�\��[y������R,�'`1��LJ���3���>3�g���2�M(F�7^u��\�����	�V��Z�>f���� ޏ�����/�fEC�zH2:=��
4��h�J��NB�D��gZ�5�-�`�T>KMay�?�N
������6[WF�<��aU%�e�dm9?.tЄ:�}�_�{�Fb�MlJ����H�1�!H��-X�ժ��a���g���!1��؞�DC߁��x���@R��T͇�lWw9�^>��M���C��!�=YV����%�����{���g�d��l��Z�=�~�䪦�c�+�Eg橙[�gnE6Q�����G?*�ԥ�"�r�D�;��.9p����VB"����`��"Y���HQ�\y �}���+Z�-r5V���� Ә�������b�	b�՜$8��-�?\V�!;�"���w�T�N�2c�̋A�=�aI^2�SU�� �3�[�k�X�5Zx6�\�'��z�b:f�]/�r�#�ZGT��S�7GAe���Gu)(Q����c��y�Jg�����L�W��!�#"�sw�4T�`��©,�� ��rUF"��;�Z�ne#���Г)��Y��|7�Ux�~<:�#Ț�ݟ"��r�wW���	s���qt�y���e��ߐ��`O�R��s�p�깪�o��&�Jz�x(�{V"��$-0D&� Η§��\��e�òc����P��m�,y�^弦����evP�`�E��)�Ns�A>م-Y�����]�@R�������Kg�-ݯ�.쿈4�'�Hk>���d`��V�2TG�P��^8����Ǳ��̙��k`��E�5��ȝ]��S�aH��]��}���8$|����'����W=��yT�; �A[\�/��gL�䍮�������Sg���yM�$�('x��rҹGX�n�|���׭�=֞i}'c��V���Τ	C�χ^3���i��>��>|9+2��)�o-X5I�	�7_��jV�b��^�K4*o�A0�W�j:�0�;j۰>%:�!�`���,�p7���Y!�
���"p�7���`L��o��z�
��2Z������&+ۂ�Q������5!=���n+	���	�'>��*��g�4����G��潌M)q�o>�e:���K�`�B�JNYbFH�=N��Ε������7wj����,h,	ϭ������Iq��X�_�8�Ѝ�iy���{�'�Y�`�G z���< ��7Α� �ٍy)��!�G�sCwoR���DR"�p>|�V�Ґ���-+ ��[���e�Ir�F!�:R���!̌�R���T՞E;1�tW��=Ԁ�<����*��&���]�\5��Ug���H�E|~N0��5�c�P���)��D�b3L�^ڠٳ/���t>��A��ʾ��fVEtB(\����m�j�ŏk�)������@����)���xwS��ɩ1D���)�1?��t)�\;�Ɩ[{|y'�	�3�=03-&����tipf�2ӌ~�g	�*�h�����?:�6�~��v��k���[��C�~H��Џ��\3��YpF]��ढ~��S����0m�&�ŝSP2ۂK%l�6�(a�A*|�+~��cè��<E�s_�F]��bv$���*��7s]+7�a��"Y���^�H!���}K��A��17� ��`�x_~@Z�X�p���	l��K8!��S_0'C,�øy� qa�Bdp�(�O.�~������8i�'(~R�/���v�g��纽)�6��������O,��m�g�-���4��[�}�3LU�O�V�	�ɓ2�?1�w[x��k&�G.�?{	gi��zP��/���@2zp�6��M�P<%3«�k�;F_�Y=�U1o�.����x��7�Yϐ������������1B�ȉL2�o������Z����V8$��a>0nO'�,�Q�(%����4"_��;%P��J����w�_�g���?����qV�W�(Dц|!9C�WvD�r� �)_ ݐ�Z~JT����=����v��q/~�j�6ӂ���,��&3�?餃y�CܓT ����ג�9J�X����e�2����]�ֲD�Rt�̻�����*�ye���8lk*WlK����a��(\��+p��?��~��.i�>3D��]��WE ��A�-RX(.� s��A��ڄ4���KeX)*�b���m.|�w]�s��d��$'��a��DOT�%<q�XlxVHYEB    fa00    1da0Й�����8�I��X1޹�H��)cDOT�M�	*��D����l�y`���>c�z#&�s�1��g3hƇ��S�������՟�ҚI@�Z��?Y�u�Hd@̱�u]g=1��&��-��W6-V��ȱ$�>r\�H}:Ǿ�o�d-Vt��L�, ?�ast���
*�S�bΎ~�h� �P"����ז�b�L��'��A��K[�}�>��o{	�#�x7����L_u<BR���5������iʜ�E	������������l�e�f+���n��W���cg8?��i�( ���x�)�s-�d�US�I�gy?ab8�f��l(���ڴ�E�n�w۲�z��l ��~��9C����uT�ǲ� o�aI`*��
���R%H�x�#ϛUAMk��0bZ�m�e(��.���y�	�O@�B�<dJt�Bw~ܜ�%<(ޞ~к�5q3q�ڷe�t{�a��f���u$��imLn]c1DW�W|e���`�|�����.��`֑�bt"�����Nz[�r��P�؈-��;E3x��y��O
5�4��JḦ������0S���u%fE) FU��S5=�_� %��x�Oo�x��Ԉ^����@�q���4��tH��Qbt��tW�U�K9>��!�P%�7��1�m�g�֒��_���o��q�^¨��BK�Y�\�Qr,���,�2��ѓ܍�G{�$\���P"�e��GM�~ǥtĐ74@r�!��hQ��e}��5%���uJ��tψW�+ۓ���j��c�ɼ���*yG��S�:�~����uƻ�,@��%-�����͌��QJ�ئ�z:L
�2.��n�$\)x�����,���P�Yvm��:���N*>�C�EOM�x�P��KT�O�j��Np���
C�W��=2����@��P�oP�̢����/ZZ�Eu�D��D)�I��\�����<��[?�I2�r��#J�򫆾eW�����7�;��e���Ds�0��	������'�z�n2�&�b����l����)�c����������,G<a8�Il�EErN.�Wlo�ee8W�`��D^�X �B�Zl)�����1��|����)�5�{C�b�m���jb������-�g�l��ݸ�!���4Mf�"�I��LU{r�gy�K��j �cڒ;7��d��8?�t����{��>���@���6v[��JXv^�y�Yw�����dؕ��7�ʟ�}�¸�~y��0�J�t��I�O�k�y��<ScE{���c����F���� �^������9���t|A�j����:��~r��+�d#B�x�,0H���p�,��<9(�'v$��A�b��� v�Sr�Ť�� eǇv��=��uS�%(����/D_���1�yz�:˱�]t��b���z�Ô�&��n&�5�.��\�ە�؇'*
�,%b�.������&s"�F��~{q�5���P���ｼk� 5�m6Ns�n�2�U��^qS͖W9�s���U3�\^���?�g��,�c�:��)���q�xk*�|[��(�^DӑM��yi�3��U�C.��o��|��Z�Ġ��k�z���m��9F�3z��|0�to���}�~r�b�$�̌���i�s|���5��w�q����GmY����B���X*����i�r��Bp���
����\�Q�?i|�w�\P��6��ҏ������
� z܂����X��2{	Kq7�㿼�����G��� o=b)�̋{g�g]��'ٜ��j�H�P��f�P`\�{�������&9��,��q����:c@_�ӹN�(����ZD�7�d�ە���1̎�& ʺ�0��ʠM/de��bWh� �3��B/mq�%~���繧�>�B�M�oG��Z�n���US53%��
���3��y�K35�'�9`��t�����	d:���aOz���$�l7mҹ��)�Q�n�P2۝�����V�}ϫ�|��v��Ʌ�"�s;^l��B��@o$����ѻ��G|�m�}��>~1	���q�,��g�7 ��yY.t�K�S�\C�q�8w����!?0�(J �'��.�4]���pm�ŏ}�1�K�Q��Ir�u�����=íC@��������CE,0Э�M�
�>9Bfc�[�yĮ��b/�a�����ճ����1�#|q�6c�,t|��zȏ�����e�OŌ<`ۼɰB��*���%Jz�f�g��N��h�щr5
�e�aE�/����&��@Io��#7	[ߥ�!�]�̝X�ӊ�;��1��\��oqA�ߧ�5��X�Ƚ��	P�:V!�؊�z!�i[�Ю�eC�8���.l�I��0����1-�̐�x/���+�.w��]�N*�!<�RчT{4�dY}JY��	zRa���)�7��"�b�Y�h��x=O_��ݱ��9��+�����Oy�M߉��Gd1����$�s��Ԯ���SU�1��MTDl4�'E�h־�J������c�w�, ���~ܨ�+�U���U4r�!nv�
��B��!�Eo��֟ӀpB�jm�sK�YW�fք�������B���O{�FJ��7^��o��6���#�Q������@�}ǅ!��hۜT��Ϫml��;9r��Ǉ��"�:����Æ��P
�s�0v��B����N|Q��g�d���k��[/� e�_�1qWW�>���Jŭ\(]�y�8o�O��Y��`��LQ��&��6���A���@E�/���P����^�����O}���[��=�2Y_�]7�*��D:AcZN��ұ��n��RL�O���w��;h�_��ďU�^���3�Q��{$\"�%k0����c�?�QM$d�� ~u��J6�t�g�I�_�g�t
:�}�P0B��s��mBD+�&��D�gɴ��b�r�b��b����VƉ K�$�
A(���t�'j�L[�t)�GO	+홟+U��s��z��3�5(�|%(�����.�M�7�HJ�����4�u�
+�>
�K��0D��������(�R5�)=~�K�����]��/@�9��?���t�g	+�E#��`����F�
�r{��2r_�]-U_�}�=)�Ų���ۑ��q�m��<����͝!�[��Ĭ|��dQlMѯ2a��L-��z#w`5z�=�b��U25�'�*[	͹���L	]��hZ&/�ϖp��-�aj�Qz/EW��{}e��=�`�*����ql ��)��řӤ�p�b3X�����[�"���~�%�H��lRB��r�.�lp>�����р|�Xɳ�5�8,]I��Z|��hF&�g��#�o����/���z`�|�~u���J���)H�������~��<jKa��[M�Zd^�0�rmʦ:�}�j�x��n����J�ڜv��t*�m��T��P�* |���vb�4��?Up�8��u������u��;H�!L=2�TË9(�߶�0GK��^��z�6|Q]�CÓ����AD�D�ԋ㪏�����M{D\)�&5Q���l஝�[�.�.�j�>�r<y��Wě�0h��b"��:.��ʖ)8EІ���,�y�B,�)�"`):�sڱD�O�q��u	�vNF Do�f�IPy���wYt]�<���d8�WL����G�N��9Z!��|g��+3��L�Xp y�Ak�:w�rm59�J/v�e���5ٗ���e%��5��ڷ�+��?H���e����fN���5��)2\$鰥���8˩�E��%�ݰ4�L�j;��{�cM���FC���|ܞ+w�_�Ԭ}}d�P����4�6K�%�e��a����t�e�L�ųdq���H^�a::��:Ecw��AV��V�e�v�̦��{"u��5U����偺��@�1p�1�V�Wd'��Qo�Ǵ��pro��)E�v�������{`�ܿ!�N�:4Ϭğ�đ��>$����6��\�K�s��l2�(����.��(������^������uĎ�m�g!:pæȹ����4j�v�h�(�%�[0�|��u^�����ć��m~�-�L��}�t�[$��8��T%1�=KM�^F�ƾrL���%;r�����[�^~DebY>�[���'-K��;��~m�@�AN'ʶ[���F�#�$����)� �1�a].�K-5-��&'q0���Rc(�v��	�V:���w�.�<$��j�ϐ�[&<��9��|a�x7b�:r�m�|�d*���}�')�N�tإ���.��łav��EX��������-K��=�u�ƙ{����,�9�A���G-�@*;\���>����\�2��J��_�~��=�)D��ǰN���S
-�#VB� ��/�e�z���$�-^��>��:����*1����^t]��1e�J�F��q D�e� ���$X�o�7@���G��l��J	y��#��Q�$��P�sź�2~�R'0H�D_��yz���|���rk�I�����m.�c&�$0ݺT@�Jδ�oٸ�Y ��2Խ�h�w�j��֔L��W����p�o3�^�1Nx�@������j�䓟���b�"$����s0�����1]<��/Kg�����b#U�|�x�I�mܱ��jwɓ�{��ъ�%�A����gen���y��G�^b��$�㉞�X��<�l�U���f��%���W�n��}_]"u\R� ("\�8?s���p��ʼ�s��]�%]Gd*X��fO��ŀ"J��O=?�ţ¾&���s��p����[��&�#�`�Q���Q�����i���b�E>^?j��޼N���Z�hI���Z�Ņg
}lc_ɝ*5�r��L�VvS�B����X�j�|dE� =��*�y�)�������et�n�g�VΔv	���r�i;-��f��wc�[���<���U����a�a�;O��V�/Opp�Y���[��|�ͶȀ�.�����)�;k� ��3BF�]��$���)�pp(f���$��w��W$��l+���{���D�y���B`�����T�� 	�f����,�����@�Y@@�Uq�"-�4�Au�=�I`�M0Sv�8'��B��{S��y$�mƒ�hY��O{������$�bL�mgT�9�ܷ�s��]�;��&f���Tw��.93�s̘��Nm1�m�`H%�>��'�ϒ�Fj�8�O8�r�hX �b����ٱ+���זk���`����K�&;,lrQ�e��$��@����p�fP�#Q�E� ���W���Kǣ(`Ŭt��C����E��B�������WZ}n���P@��WB�KY�E�$�}��r�D4e��}�v�v�#V���^6kX�����Pl�u4�릀t}��=΃R��)0%�cuΑ��p�q����e�Bh�Ң��K�V͛���$XmH��m��:H���`�ǎ�a�����t���s�V'-E�)��ɝ����`�x"�%/Q �Q��<�/n�L(��Ǜ@�y59?3�%��	����a�Bx8eJ�U�i�5������:�1g6�^�=��T��� ɠ$�w�I͟�%Ǹ�V�F&�{����QTi"Q�Cy���~Ņ�a>��j;���.��ܴJ����u:Չ0m��c؈M��eSD�C�T-��s pמ�	��u�I�<�]Ƈ�:j�0B�ϊ��ƞ��(��rkf*��"~ ��!tv%�Íg
�ǌɻ�JVWX�`��"F������>R�&��¹��(�1��?S�����ƌ���<cVZ���	k#�붼6Y�@2�G�9�г#�2��)����%��):�$ �ϫ�,eWIl\�-�$�����귴<Jygmx��,V���j�"��$�"&�'�DO�`���;K�8��c��-���k+��9��pe�^�,b;���AT�'�y����;�<��[���ޏK�zlETH�~ld�,d�.�o<��P�_^�Ū��xv���!F�BѕZ�,G׺�,�~-JG����FA�\N�ԟ��]΀L��f�NT}�R��_>�ۉ�?����ؙWa�l�4{��Ep��4��3�c�'����a�$C�3�D��E��ƚ:���b��QM��uf0�6�^8	�I�0�,M�]c������_���ʪ��@A�jj�y����J,��(�x創:*=ʍ~��T��,a�G��zv1E	��tzʮf̫����A�|^L��<�J\[�*��A�{��$@>��Q|$0 McG�őh�_3���
��ͻn�S��'�2��5tXЂam��i$cw���6��[J�a�A���z��.Pb>��>~a�CR"�?UU�sAN�'��#7g�Xܦ�8��Z;�2m�3�e�X9g�@���S��S,�B8���#2����3>��Q�i�$5�+�e(�8%1���2�N���㋁1������CY�_8�I�=�ޛu/�EU�\ݚJ'f�{$@��l�O�E���0��u�v���|�c��e�C�E(�;lH�}X_	iN��� uJ�8PGS�;M���CwoH��w��I�'�E4}�5�Df!�� ?�n��U?����I/Km$�&���Z��,f��X��P��菲�>~�|Ǉ�ICo�o:�;;�Rl�����r<��%s��w*��Q	B	��v�o2V�b%3°�3�	ዞ��8`9��q�y�>�Ј7���e���G�}HM��_�WEL%�i���É	���tf�n�=�aSjU��b��{om�7��Dy�e�莴��d/�^>E}�����,Á���(g��*�����*��~u�4T���0��=(��ɀ
C��d�G,Q<�;�#�5���B�Q�R,��8�S�N�g�m��V�Y�a")K��7�]��|uU�+�,���(4/�ia�����
�g�n��AF5�C��X��/
�kq��2�/��]p�
�������^i]]���Hn�ݫ�\��?IO�E>�T ��B�,�]F�����/�;|��H���*��B]Q!⪍��P���I10����6̜���Pc{���L��L��ɦ�[�u�#$�f-6��|��??�{r����
��%��u��(����hZuϝ�`�/�~xC��΀�E�v� �t��.pyZ���Ə,Z�u/��T���{��p�>�W���B?�p8��-�͜�7�{ӱW���6���J'�����?�j$�kw=9����(�����I�B��b-��U�c)�}�%{���&`zK��F������ DFfG��2ݐ{|C�/�������|*@̝���7����y���p����ț5므<�-�g� �ev�*c��R��� �7c~fZ���ȋU�Q�7�x���t�95�}��9
�b&&颅��pP�w/�yD�Nx��l���yx���A�:�pe��z:Q���U���y�IZؙ䟤z��&Z�Z��<O�o�9mӡ�k�C���H���d�_�n���<&�j�4��[�XlxVHYEB    f314    1b50AQ�FQ�4iv����l/�:��d[�;
�}&�A�9� �2�A?}q��T!�ڂ�#� �L�1����!:�O��L���N;��"K?^�^J Y#��}�/h|]i�2P k���  ����:sF�EM�x�ġ�N��x=j����BL�.nE�6V�[���i��˯ܢi�e�!�(���5J	!��V4�Hz�PY���k�R�:ҡH���um�\RP�v�L�'�an'�2�2r��F�������>Yff��T�&:X��<1ղ��?��
A5�Qy+�T��ʒ%�YǹrJ��b_GX�ֻ��Kd�
�=e�?��'H���-�����6w������f��mW�y��_&�����K�Т���T���.qE�[�:��?ߊ��?�<Q+��[���轲74�LhF�K/Z�sqgɼ��3W�'���t-��:���lz�S.���x�{��������ij8B�oT�����զ��Pv�I�y��#�P|�1��ۄH����;Җ��~��{Hu}���Y�6ҙ����EM�
�Գ�W!��˥S�k�ݝ�zB�.O�i}���j��;��h�4Q�M��&��ƴ7B�j�u��|����[���N:���-��g�\Zz(R.R
��l�Z��.$��YV'&{�?j�	��f�L����j��55)aǮ���jN(�F�{hԛ�9��vL�yY���)�JE�QL�-b0�q�]��m��by�_�Z�l���7��x���VZ(zS?�} �F���n]�kvz#L����5>W�;�.%:���S��W �p��c��n�R{� �'���A

c��@c?lk�'��I����Q'o޵��Q��,|�-�y7��lӨAi�t�X��R����.{����ْ��꒟#�-�O��O_�g�
Pi��V�5����{ȏ�����N��h�$��߽��9�:�����36#P2_}�Q���?�Nt�bs9K���c(�gO�(�8���>:%P�4t���$���	��{Y�nd�_�ԖI�4R�Vb��oS�+�|:��!�bLG�#�u(F?`'v姽@��E?�]n�ɝ���6����� �w~�%��м�9D9U�� XE6S$;���e`�$�_GO�d��T�R�_Z�0�h�M�j|b�����d5오X�_�HGU�p����X
_%u�J�5����>р{���_��=WQI�n&�`G&��a��H���������2 �Q���ۊ0��Z�FT(�
����B�s t�{N��v�9�R`S���k��#p�E���ǒoR��$&�G�0�)��+��4H�������f��E����2�
P���M�Yu �.q�M�o�fˤ�P�a4A?�^�Hß�}�-�l�q��C ���4��)��D��4����*a:��?����*��UgL'��TV����+�e�5'U��(n8�a��9^M}��2��,�Iu�K= C���>W�k�* 2";�C�ע���7M��8�R������8��0��E�1�*�(mY�7A���/ߨ嵧�2�Lg��jx����Bz7�Wn�3�yz��Ph��\s�t�̻A��)�t5BbJ�x�x�|����Q����t���l!��Ҹ 	q(�Z�ʱh�9��ϙ��>���_�I���Qp`�Vc9�M|�E��m#���(Z�,�]la�/���[>�uS��V��~A7��3d���Y;�.�p����"�-ѩ��l��[�}���l���ā~/Xoe�����;&g?�� ���nm[�V�'1F��������t�j2�;*e�������� /��H�t����2��y/��oe]dj	-"����}BjP�Tek�p����� }f�ޭ�qc���)U2��l��4�����T֧�����w��|��\M28ˈD����X�ë�/�v�~����}J��C��Pho?X�����ʹ��L���8�4�x�|qݪ\4�A���f��3j^�*�t�hV�8^�M�dل
�uA:
a�� ��/)DL�ʯj�x�t� YȆ0��6B�����`�Җ��u��YL�~�z:��q�fsB\c�J����p3A���M!T?	��ý��j1�
�\~o�����"����E�񂻦ݭ2�Z+��c -�عP�q�QBZϼ�l�m"Sp�wѠ��@Lk�Ā�s��ݽ_�c��̈́�A�0ĸ@��le����;H��O!�S���c���Qc��b����i�|o(f�+$[Z�2f���	
z��0�;�K_��G8uDAO��Qc_�Dx>�jl|�v������o��W�^@oi���f ��g��y6���B�uz�:~�,����Pd���P����Xra-��M���aU����>r_��j�m�1��R�$:J�^ ���AC�h�P�w�gi�3�n\�(��d�Q�� ��xL�וֹ�ȕ�:�EP�u�<إ���1�瘔�j`n��H�|In~��U$p�ȅ���<k�
���ɷ�McA�z�Wl��`eK?�YL��G�
+E$�9eԖ;w�5ᩞ>� &F�>hX�]DC����`�$:���.
���Mb߃�L
1C��򤝧�	���bٺF�s[=�4��\��O"�O�\�b���^s�@�o8�J�i7���ah�0��P�T���W�(\7���y̼	3R{��L�Ȯ�MYD�,�ހVG��/�p��B*a��.�����i�wK�!ͻe_y�b_M��*�l��<��0�3#���GR|/���5��sQqAA>⌘[�'j�L9�o�njG����'��$�҂���*�Z8��|1�![)�����ı�*O5h�Q�ے��Q�[{��+�������M;H�!���hA����2��!��qc�JĒ&�����/���u�7V�hPW�r�S�;>*|t��B{|G����E���/F,�q�W��ÿM`�R��5���͚���>%> �=��F�H��c&� �=�t 6u��LwD���WxCU�(�'7
��s�]Z���[q׉+9@���w�3�h1#l+ˎ?%L6i�{&("2����j�3�Q�_&�H�N�: )9�:�Q��dh(KBY�G�� �5�V�?��ro��#�S�Ep�"���e�7�~���� q;��L�4�׽��S�_��m� �+��vS@�8T>Z��d�UJa+˨��h��?�����`E��#���#�1��I
�*�~$�\ѧ�P
Lq��uʐ�������s,�.���XƚC��XZ��lN� ��'����y���WY����KV��0���k�h�#�2� ����W�/se�(a�ac��O����`B�Jx���4^!4C�\<&�{M)U��\��5��o�8϶"�v�ʁzR��SVݟ��*/.��Ŗ-��C�/�w��3@���t���,U�l@��'��0sgh���Y�"C91#lT\��B���`��2�U�^|�%2%�HA�#aE<=�g�#���£��vtS�5o\5�frѽ��F��l�����E�2�׮��,�����A��>�}�Dk�vj���ӻ�S��_�OL�M9[|[���Z���hߵ��
��
����0��?�YL�pƲ)ܒ��A�5����K��;��q
�Jw�;Y��O@Dj�
?���Uu5���>���B����(��5��T�M"ȳZ���Ԛf�N�PYu�"�4�e? �"�8k+����>B��eʆ�;�cu�T�O�n��`�L�+��^�4�oL�=t����u�1i�J�m�F��	T��+-/#"��@��_W�6�D���{�E��{��?O��~�e;�Aga�k7�GӧS�#X�ur�+T[̟�􉨽tҢ���L�e����F(η��V7܀�����ع����a�-mR���KZ>ZD��+����ã������ѱ=O���9�+x��A0J������p24���qT2�IA �d�u�̆X�������3~���؇T��u���Xe�w����6�R�w�I��uע��9о�~�$-[v�H��K�'���&���OL
aN[3�V������쥼(����11eAK���,���O�lE��m�Z�>�\����T_�J��AᘯX]��<,(�ČW7@�3I��)��.[�"1z~P̓l�n�[vT}���e$��U��NQ7�yQCR?>�b6���]�u�IY�}k��l)遢q;'>�`T_e�&��g�l��	�C��a�����%�~ĝ!�tr~�I�RϥƲ0�po��&�Pe�H�a����UI➜�B��u����Ss�����U�e#�U��b��k��@��K�~`�MTD.f˵g_��9�=G���F6�X��B�����Q2��ēvqmJ�2ʙ��3/Y�Z��s�>WI�ޠ�.{�����mE]�{Ü���L�G�J�?�$RM�7+A6/N"�1�Ɋ�ʎ�vp����� �"s$dD�]�»?r��0�4��RF+y�s�BvҴ��^�>|p6{~�c����sX\ms�1�Q���n!�I8�%+٥%糉�.��\>��bY��H��8�����qy&F��1����}�����WH�?F�1��xԇ�֑6�달�O#$��び�h��p�tb��֩��W�b�@2�	P����Y$Ș����h��]�	���\���6w~�c�g�13ɘ�0��It�Ze�1�H=�є����+���@���ῢ]���Ÿ�ޣ��&����+B�0��P�J �|�c�e}9�������E�S�U.̱���f���/P�5�w�t
�Ȧ�J�m�Ď�����\�N�3̠���J��f�D_�z��mI��Y�n6���ti�i�;�����0ns�Ma:��KQ%��������Ͷ�ei�,h����a��:\c�ᓏ��Or)��4���t5d�@F.G�YE��Z<�|5(_R�	�;�L��'|���PJ�պ>3 �FI�E`{� ��Q�QB�[e�H�&�)G��?�t\��kyY�p[C�������`0�7��>�����Z���&�֙�:��)���3b�}����z���d:������� u1�=����iyp/����64��C��?��hm�D��!�P�,Z߳N��q%N�ԩ���D�p$�ϰh�	��#���{*[���Y�����yD'p&UmNN�uy����ε-;�Ubā�_x�0��l��fy������p-@���7�jA����-1|�Ie-L+��)d*(�_�C:T�k[<K��lS���lwD��	��]�yi�;y�
���Q���mU;[I����K�sz��E0!�ূP�d|�}�4�˜A�uiS]�}�<tpI�Nܸ?"t��k7o���*�V�X�"�q��j)��b-j��D-͡2k-����X����sb����B�4hd;��#�|��#F�H���E&L�p}d��֧�yO�6j�umZ[�w�����,brc=��������mj�P�äX3l(a'D@KJ�{}���{,'� �iv�s�Bೂ�đ�z�X[^�z-d���b:�k���|�>%=���?�a��q2�$F����=�f� #,�:�uϴ���y��[�^@zh!]�-�����A<��:��9�o��Zh� �-�9�`e�~V��b��I�;�c�Q(� �Y��+]	������o>�dh�L�M6����O݉�T��0�Zs���y�D�<2��pV�����R'u�����ǲ���6��iAE��hg�Y���uoA�٥�-��D�j"�-�!�$BQE����#���4�&%.�D���dp���0{�����=��y% �Pآ 2��9�GJ����n����h��2	>0"NS/��ʿL��b�G�p\�⫋��_(qS,����!��SՑa�n�;��f�!1�Bk�]�u1�T,�T�A�� D�����\��d�Q ���cb/hF�YҌ��1 TmnW�Y�q��h����q�>{�$f�,�I_šGcC
$Zq�q5��T��b��%�k��FU��f��9�M�ħ��ݕߑF|�A����<<m�-QC��8q Kx���ۼ8"qHv�֢@��D�"S�m��6kaC�)�X$.װ8YBk�B�8à&���"����=}�
L=��c������U�|�ⶩ�e����V�Rڥ��m��Rcb�9Ĝ��iN�)X/#�>:��L^��x�Q_UB�й�X6���lD��J�����ڳe<��O���*	���D1	�C�j���P��+����5d�
a����kg&d��7�d��'[{���]��}x'��q�#706��8?7���Q�lzN��C,���Xoq���,)�~��@�kz%pP%��� ��a����>���rp3��(�1��,�[�{V�	��J'^"��9hs��^�z�)��+�k�\������N�_U~+�6��>�����ry�M���$/6�c�(.��ޜ)L�O��: \���އ\ו�YǪ�0Dq*&��N�p�P�ly��EzebD�N�V����D ���H��=}�r�k���%����E"<YӉo�q'uDX]�$���c8��{�p/�r����<|m:򳮐�|i1��u���(3��旾�!q�����U4�^�׼%f��S����;.ЎV
�����5�����A��V�&���z=�R�2�:�ñ� m�4�0�cL�]$}�'�q��=����	_x�&P�_�M�e����nd�w�.V���7N��`��9l=J�Q��Jʕ�H�.|O)�pC�gP�\󯭑iw�t�x���X �����U�l�S�SQ�M?Z�����ä"������V�tب�M3�%��q�n��{ߖG$.�����j�{3x�'+�3h���W+�]�(���fb�2:eð���m