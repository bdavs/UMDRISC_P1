XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����*��o���d=�[�?�}rX���	���L��@�n�Q$(]ܢ+h������S}JQ'nе�A��B��N���p�78�LcK&e�Gf��5a�z)��`�=z�)�����.�K�F�ùCo��{�ϞdIcC f̍&���r
�},� 2
pg�J�-活AW�9C��ބv���Ц�h!.u�/��n��X�+9��MJP@�~�4ғ�M��vl֢B����y�PȢ���h�ia3�7��vԞ��Nv�bU0����͐�4;�y�J����S����Q��a���� ��r��*�m�1.´6wQpo�1&��­�wx���`����o����j�͗`�#�Y�P@]]>�ы�U$�g�?@ߛ�>�O�*�O��&ؐ �K���"t�PCut�bZ�x"�wX�-�נ����5~HaT0FDO{�D�pz�l��6����7�OMq�/L	�� ��ǭjw��'grŔ꾙�؆#����-��zdI�B��\"�cm�7-^$�=����m��s���$L�V;��Y$��a˜��?�@��-<h�6�f #�Z�P_��8�^�#�6��1Y�)`}�w�J6�����d�\h)�Y�r:8;�$ӹo��`V��eU�O���`�i�ޫX�q����?J��d��D4�Z�g[��.62��n�;���{pS���;��4��ख़I��UZ���E�=���F�V�"�w��{��x�b���6��}�ڮ ���M��A�.s���pv�`�7/��8XlxVHYEB    3042     c80�\"�@���U�J�F��q�T���R*�T�����(�?�1�O�	/�iʃ�2���&�E�Lѓ�
��E4���$��L�웆����'�,@S�<Z�ՆQXe)sn<�~\�]�b4�!!1y<�>7ڑ��D[W���]�?qc���V�ˀ��H�KW��s㡗4�����\�/�Ǽ��`�4�_4�b7��~1̂�h#�$�A��%xK\>U�N$����7:h���"����a����?��K��}�*l,�߉�O�4R���w��[�b2��.p���u�Z�W�|��/B/�a�N�*T���:(w�8�)O�ȬJ�#���d��p�m�Gb�NM���"	'�'ql�PF��Ӗ�6��2z����%l��cV����x=R�!x�w�A�~��e�0�r���}>Nk8�"V��t�j���wu���P35jw���l�&)�7b��j{������A��^�ݕ�u�w���]���.��,�BP��	�6
X/�=�s�ZWW���Iw'����	֐�u���2k��W`>�?"{�gj	[n�G�����p��i����H�v�4@b�`��y��w��_�x�7��g��Ȱ�'�rҷm���ʲ��&n"H�b2n���v��A�0溢�]顤�E��l� ��u����n�G�������(�}��	�@�B|�4�b�pu��}+)_7hʴ�'-�.�-UO���ү��$��b4�=��ö�K�<'5#jq��P)�D�6�ſH;��7T�N׵|Ud�ҁY.�1����gF7�Z�M����L�h�D�ο��L����ϑ�s��1u����x�XTo9;���H��=��ʬ�հ�|�@�s4����1���/x��ٮ�]��*�#ӵ�s����Ҝ,s�<�*�~�v-��FZBٕ��$���Tһ`�s�� �@�p�_�+݋������>�(��~L��<�cmAU�=�f��cd�hf�����̰��wǡ��H�}{��ɐ̒��s,��?U��양g�hh�p������M��vp��x
�(n�GOW ®�a؆�p��Q{(r�z�v�^�{'���Bi2a|X��O"�G�#2��֖_���N�L'� $�R�g �4$�ZQ�+i�z<F���4��`�+��)'^׻���P���*�Lsk% #�u���m��n�����˲�_�����{J�_QS���k�� �mu���,�!d�Q�96��.���b�n��z�ć���!��<P
������p�� UV�)_� %�<N�j��_C��x���J���ҧϗ�� �f#]@Z���Κ����hQ��`��7^�Nq��
�,�b�Ζ�K�e�ݗ൮J����ϻh����=ݕ���;VBA�ϳ��Ť�l��dX\c�Q27��1���--^E��R޳i��)�@]c	�(Ӵ�ݐ���<��o��:�L6�'��r��8u��<�	�7�d���)q��6)��g5���zm���[�2�}C��_Օ���iN"H����^�&�p$�Ϫ�Jtį �27���燘�r�X"h�F�=�BPXn%=<�eV��B�l�]\��׸֗e���b6[�"ʃ*��L,���D�m����X���t��9���OǾw/U�	��'�u�5�ӟ�`�*�3��N����e��#��@P�/�]X��A7[��%��/��$�W�c�F���+�L�"4�RiO�Cy/���
�^�%Uk��(�-x~e([�O��f�B�I�W���Ќ�ࠃK���0(W�&X�\�d�Gx8��/��t<3l�j�j�b�Ba70�(!0�C�%_+lI��Y�hR6hY�/�Ӛz����ߩ�#��݋(p2r�WboVo#��mX�q���4-���m�9���#�������k��EH~ �Y�]9�f��Ny�'Ő���S�Z�.j	�l���d�x^� 7��S�*@��j)b#.�澞fb�q;�'Q����)�Sf+��H�aI�}
������G?�	��qA��`}vtȩI��Q�~v�,3���hRt�y�\�Cz�m��25�]� ���+SE�-��� q�����G��~����[�{��v�ʔ��&���y��.[@��Z�L�sZ]�]�q�)A֋oڸEW�y	=i*��B�
v�ta=A�?�\L���N�����(��5c��5�!��T��F߄����A��o��D*ri�&�9c��,�BŪ'��9��C�͒�1�W^���@����xFQ=���uVl���K��*T*t��Я� r����gN����d?��oe�r���7�;��7�Ԕ-j��GQ� ��	�����|*v�#¿�]Q�EG���Ǩ�v�?�<H̼l˥�3��t�Wc�G�"���7��	�&6z��%\����P{	��Ƒ���B��q��j�>ܕV��ⓛ(�����w,�O&����f$��_�Tk���۵�m��2����p�>H�)�����!$�ܗ%\�,��,����σ$B��#����w��o���}���cI��'�	c|"O1��N*�sL�9�&�SF�Z���>��`�i}L�㓹An}�iF�9
��h�̯
kJ�Ҭ|&+M�K�9i\�ǂ0��@QT�+͒��
;C�/��n�Э{���j�
}�7�9�/�P�x,#�#�!��|��~�H�ɠ�,�St?)�۸P,�"W`�]���l��1LY�=@�
�{�?����HF0;Gu��u�U��.Qd����Ӝ<�-��o鯡�.��8�Wc��xL�|���U�o�yC]<	b���
�S���Z��FF��i=f@�WO�<��K����p�19�U����dQ��$+˔�o��T����pC��=sH|�l���z��܇�!/ȫ�!U�j��2=�ؤ7�>�����`��ȕ��"	�TӍ�bGu->��W���l
��j�l���)h��`h&ぁ�����k�?��<�iJ��.U��ܯ�6ޕ �Yi?~�x,HB��\+�c��>v�I�y��ydh��.e�g�O�h�t�Nj�bI���p�"g��4��G�9��=�G��k�}���}����Zy���YDD�?��}��*h1U