XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���qI��М�0�\�p�Ԡ�Ըx�=�08D��ګ�J�_ίt��3��a_���|\��� ��C�PA�!�Hra�o�'��(�4�7i����3��b�h-H�;"j�g[Qh�}��o�:��Z���V�U��8ڑ%�R��t�C]}2�L��jT{D��
I���;Nd���O��E,��Y��:"sB��:���N���%����g��Ծ�V�Y�o�5��+Ӄ.@T�z0Vi���R�~��p�v�H���V������;:Zӝ{!����R����䡝&'1�¢����M�km��{1ry�m0�];�zh�q�T������[y,�<�0͗T]�}[n�*b]�,�����F%��VS-=�{��������=����R�N~��P���p᢯V�-�p󧪢��{g�TԪ	�۩@�y�Gߏ�x�e��)��1ݸ��#@��42T%&ΩC��
�{g���6�z�O#.�v�� �E�lovf���}���ػ8��9��#-��Up ��9le;�'��a����9�l�^X�
}����r���㢓�!�.��s|F�e9����f�;h@�>+Rlv�Tl���
d��&�/�~�0�s������(2�uڢKL2�6'� �To��d˯��C��A�4�>��בn�(V�P>"G�����u�)B�16��*ࠚ�!u�̔l��U�L���2�u�1��.�V��QT�G�C�<	KuX���.ûo����8Gm���DXlxVHYEB    fa00    2910N�*��AK��+�,�䶮����W�ڡ`�����΋~��w��fB�|}�3�x�[��#�����mS�iXP�j
�a7��vw�|Cb"�ه��$�y��Ǳ�{s�~��"������=���.0���QnH��B��,�"�=7�'��4�GyY<���\�w�&AVi.���)���?���>rsaB�$O�2���� ��($���Ġ���7�grq)��s'�w��PT
JW��!�C��L��):a��Jְ���E�D �W}�y�1sR��,2��D�Oۛ�VX�=�wO�^�E�B<I�����_�5u]FD���hC��� �*���� ��]U��@0?t��V%逿��1��t���D�Γg	��iI��Q���#s-�3�v͢���/9��i<#�`G�?���o�����6,y�;�`遍�6H#j�?�|vB��O|V���aX�W�@�ܡ�Z�Y�6A#."�by���7�t������.�ua���tZ��c5��=@$��M�v�=�?,����n)m��w��ЏA}~p,�s�]䄢1N��Ph���WюQ
]~.�']NgSA�8�1_��	኎)���t�m�����j�i]Ȟ	guǾġ��t�O�)��} ���MI�c�Iv�EeQ�^�^fĶ'� �w�ΰ�G�w���s9�vV������6�&�Q���f)W���@B���[�x44���*A�Q�r@},��\C��Y9�e�Z[��q��r�z�n:vw�����Ƹ5۟��J��G��C�/��6��|Ҍ���xXU��5Z��/ӫA��r�t}^�C��%ڥk	���1Ͱl��B�t��+,2{�~p�R�E�d�48bNd�mW,����q���HN�WU�/v���cn�b˲_G]C�
�hgڂ��y;`2HO¶�Y���H�AZ��_�y�pC������
��UI�gdKu?
C�5��y8uC�%��}��(}�4��x�-''�}�B�rgh:S����q�h�<����"rU��y���Ȑ��S�rW?{����?��/p��D�Fj۽r�bCt5�(E5$^M$|L��pw�D1�Ǟ�L�]��ԙ�+-X�>�a�c��J�0ni$B�@���ʟ��F���y�2c4\���*�!���m.e�mz��&���!~��2�I�5�Wn"MN�o��V�̲��<��s��}3�g��{H��Y�0��.�_;�����L��j�vN���>��A�;_&���U������ l������%$m��k�v�n�G�A�v��G���ϯ"��'��2��Q�-�u/�WDm-�?**�W���c���,��:1Y�f���!���
��*��%�F�$�?�`H�_��o��{�N�#'7���+
��C�2q�L�:�T1s��&�0�M��ˏ��tFM���4.�+��Ø�g[�h���f�&ld:���'c��oS���BD��Kp�8,P�q �c�K��!P=������G(�9s������Wt����B5u14@ �����?����	U:�ָVxL�����C��~�+e�B���.��,S'v�Uhkq?xYe����sƏX��5&����n�t�*����;cJz�*^ѵ+f�v��#�.,�3���Mvl�r�n͈h���{Љ�o�GB��W~+c����A�F(.�붞��RH:F 
`��qL�t�?�{��NB;L%���=��1q�oj1Yvb��pe�i�����+x�	�Z�6�g@�g��ڽ�ë�*K�@i��!ô�	�����G�!�xK&��璒XjX�-�����˰mӷ&���^��CÓ�0Е�ퟧ�,�hV�ڞ��T]�0Y��q����=?#fl��O�{���*�e=Z�2� 6��j��~12��:��X7��/\��W��`��aWa�
MgM[r�~����u�.��֑hi���ͪ^,��ڒ� x��踱��r6,�,����'���e��EK�hu>�S~�LAj�'i�.���-�x�?���vT�|�<�{�#��oYhi�L�|�?sX���H��k� ?�<�wן�Lg*����7m>�����cV�Q�iC�x�}�>E���;��SSܹ`I�,�mXr�׎�$w�OHQ/��@ao"���j��1ϟ"�ROD\m�~�,tl�Fq@_�F��=	���F�&[x���䝆0�t,7��Bf�ٮ*g}CP��ovvC��[�L:UAQ&�kk?J�#�B��?��M�mku2�Su���Idy)��J3�����4cu�~�+B���u�Ǿ?���v���2FJc������rp�m�ɯ�Brw?��+������^��i>��l8LJ�D�똚�6VC#Wq��1��LGr7��ĞʨxFwX�h�j��@��sO�B	�o�99��1�+�u���q��?�~����r:���/;����#��:p��<3�
2����}������7��~]�(��f���	��$�M�u5 �@�M$�pؓ�@��T�i����x���QX��W9Gwž� "��(�	����p9Ǣ��CQ�-�sv��˚�>QR~�.������f�8mյ�����x�@���z��k�/�>�VV�%�*���M^�H�e���0:�����͑!�y��|J�,�GF������������3*�; :��W���&� S�+%���޽�BB���!��T�ʸo�
��n�pt]v9Q��'X���w�zYU�3���^�J����=E1*�g,(Ghy�X���F/�[uXr�%?Z�<��e�̀��G1��{_2<ڦ��q蚷�s����N�4Wݸ�2̟�&�`�R7�u�r3�K�2P�*w}���E�;,�8���s�=&z�k�:1p0뱃8���V5!�NY8���?HCu�=��`P␒�7^�= �������#]��/|PX���������|��7g"�_�oP֚n�E܁&��V7�5����������@�Ԫ}��N�F�]�\�U�3��%���v��ye�R��dq����2�|�O'�F~|~�����c�b���w�\tu@�(0qt�����j��Ss�~�|�"����E���J��/��b8�-���&��kW�>y��R¨��\�/ph�R_��'�>�(��twg0�>���C�_��O���� �P�3��M�r��QZ�߇�
�x����������2�BX��쨅�=�p�4�����ɿ0���.�l�7��/�2���2Mw��Gws��W���h�@�f
d����d9�@KO�R��F~�����P���qv0T�S��G%g�N�}�Q.�u��了Fץ���(�Hp��`�gsl���	��詜�C�E*�g1������������ˋ���o����Z}�Z��ɑ����X���qSd�M8Uw�A���Ƈg�mj_�^��:�o4O7�&��6�ԋ ����Wڶ���n F:.���^��B�W�o�7q��n1��s1ۃ�9�Ŗi���{L�Sb��x��,\�Zmc���J��Q��j�Z���J��Z� bAy��OP�I��Ņ�]�k���w}��ş�6��ݙ��B�[ݺ�i�3~^�ݣ��L��*��㧸��<���Q�ɓ��K �"�K�w�u?�%�������m��ͧ�X����N�������0��f�YRs�fK%�-���'	4��a�S�ɾ@�2��c�Xm���ћsR� ���r������_@���6���s���j���H6��4���}�c�U�yL�Nz������p�i&�3]q��{�:����QeK�����K����R�&�������>9qt����ٴՕ.�p�a�[}7M���=��V�_�?0a��"QB�nu��X�G_��M,�\��<P��2��scx��z���L�_�Y�~�tȬ^d���6Sg��K����C�xRr�cy�Iw�>�_W�,0&7�Q&<��Z�0�a��"�M��;���K\�Д.pX��F�P@��(�.�7��{�����U�������Mϳ��̬�l�w9p�����v��1s�i��z�F����ب[��c��d�͛��/?���cg�>�ݯ��>��~|�4�T����F�Q\?����-���
����s;��d�V3~��n4�t�s������ �
S�( ���z�D�3aH�.7y����I伧�N^)�~8��^+#�IjXF#c�U��9�6����A)��H����cW� }B�#;�^>�?���-��b痴T4M��g+�?Ub]E�4�ˈ$Cf'�]|�j�-"��� )W�l�hD��Y�wU=/���0~bb��6.J��[܂*�)���<WP���@�4�L�D���hϭ��������'oƜRƔ���T�x�Nj�0��{_��j@��t{����M����(`������É�=�N'PS�'{��"��7�D|EqH�b�oS#�ueղ#B��/��K�� >�2[g����y�����:���:�0T*�޲>2�{#��!�Lu�/̗7m�x`�K'�9�����S��\�55�֩�3����`�������^���KBH�������G�OПBP{6l�GҠnJ�%h�� ���f�vo����nR���K;�#��p!?8���~�Q�V4hk$<U��/���?��Ѝ0Åʏ��؏��T͹8�X�xMș�0V5�=�������W�b����ೃ��u�:K-ޖ���<�w(j��g����G���Պ�(%'���`a4�{�4�J����<y5WP��u!�L˂�L�,��R��Zlb��~��h��4�`��z�<�x�+��p[h�݃'ؓ"���!�S����u�������������D��ե滫���E6$/�&�{���{$�|�[xyLZ�����ڂ�ǧ���;7"Ϩ�'6�.�	�w�/�m��mY�J������dOP��˥@���]���	Ӄ0��3���qHvB�ES�sl3鴋|���1��<�Gى3��"�8�:�L�ڙ�NM���ET9� �sr��$�"�冢�]�K"�x���n�}��M�Ǹ�0�=��΍п:�.�,�!SR� ��$�u�TB	�gYR �� +z�{�_��܊Q%0�__堸���~xF��r��n��Q�2>��(8&`:�{ ��h���E�M��@�d`�9+X��I��Lʸ��ّ�}��Ӑ�[��u���f�Rrj�;Q�Z���dZp��������Ջjm'"�y�;��L��k�+�"��pJY��rk������u�j_�����z�)k��a�NO������!���.�qïEn"�g�U���/[�@J�#��w,��L�	5�c��T���(��(7K<��� ��N �Z��y�2�{�B%���:.1���"��ˢF8�Z/N�Y��^)��c(b�� �Rw�h���giR#����Xm���۪��!�ع��\Q��@��1m���Z�g��\�(*T��h1�&���ʫ�sAB�����_N����#i�~z�X�e���F��6kA���G�7O��S ZS��,����;\�K���Ua��m�į�����1mԪ���Ê��_uU��:��5�yPN�4��xHeVݲ��k/Mp�4~��馳��~��/bT�ȱГV��<ϭB9of�����_D��-$�ZY�{�	Y�*:�w���K��N��x�s���hgݭ�{�83Az����t��է%��0P���}rԾ����y�1��3]8l���-�ٚR�B,�	9#����~����Z�//!3��M������ܜ�*P���q"/C�9�+iM�M'��n9 ���j������S�������b���Zqy�����a�e�$w��R>>�tQ���T����v�d#��5L�����{v��L��8U�F&�J�r�R��J�U� Epw�0�Pq|��h��J�8���$�9��+�h�l޻-X:� AZ��$r�@c�)�i"I�[O��g2Y����=ی�C(q�<��%�n�|�WTg/m�b�O�5D_mȗ�jR�ߐkuVzE��l�R��ˢ���t��Rfޤ���˜4u?�Yֱm/$H���bǪf��B֠~��iN����]����:z 닿{ބ%�Q9Yh��	����n��z���#[���"�u���">�
�d��E�G{�E���ҁ~�ۈ5_��U��ռ~�6C�HE9��.��g-O�������L�{F�@3��v�#�TW�5��LY��%�i&�Jr��o�X�**tk5d�ae;�$�ы-	�(� Pן]c(�M�n��(��n��t`ߺ���~Y����4�e����|��}d��.���I@g3s�?|]�Nc��hת�B�S���5���'��>���]���V<����=����au+��C|M^L��ǲ�z�s�4%�֒J� GQ����C�c�1����~=�M���c�ϸ�$��
��K�Ø҅�������cme�3H��6�HXMƷ��;1܁�J��^�,��QG��<�o�+����$��x��z��OP0Kx1rRa��Ȱ����� sM�ƚ������?��p�PC�[�x�-Ȏ5��~�;�lh������,���d �Aʝ���c%P꿻����$��o�⿞�W��A�>�'g��x(�4�}A������n�r���G�d��d�@���f?æx#s/�eUz�f]�=�H�Ĉ�?�e��3a ��"���I �$WtmRGK �2+k�Kic��m:L�{� N8�._�K+��:�X�͎1�4	R$�%^�G��Łt�!�-Bt��3[�����)�����P����j�pMb�������ED� 0�"O�����f/�[�V�}�@�������.��{wL�Gw�X�[;�]�7~����e.�T�5��y�M���9|iޣE�N�J��9��=�(��,0�b/ԨG�S".� 
�0��Zη�k�}�qʍ�r�ͫApT�!ݱ&n���sY�"K��C �����A��w.����gO<3J0���{ӯ$qT�E�p�7�=\���J&~��ȝ�@�Q�H�Bݿ���h���K�
�Y����\�ͣ��s�͌�r�|y��[�V�l1{�����\�C㏔G��l�a1o�kϟ�\6�X�,eW��׿#����jQ�3��^��~�bo���W���D,�Wi�V#����]��k��n �����mY#U�*�b]	�HY���f&�������90U�Z����)���hf�>M�^�r��?����ge7��>r�Q�t��_|<@�/a�4����m�Q%�BӼ��B杻�2�0F�O��0?D�m{�&d���/��b7|$���� �6&(�r5�����O���Y��� �^" Y�B�h�-.\B�:��Ap�>#�7sV|�>��5���e�BG_�-ށ9��>���Y��R�A�gD�|�r���ئ?i��:1����i3i����W@T(Ԫ��'M��*�$;b��x�@�Q�Y��Pcg�m2UQ�Bo�.==��q��܍���2�t�"4Dv��A��|t��H���^
 a �=>)�; ��^e���	"�����\�'r�O�n���#���K���t�"<�WT%V9Wo>�1��og��j�(ep��0LL�zX�~;�ǆ�;h�m�Q^bH���ǔƯ�������bB("j`���X���h��]C������}����K'��X�����ة��;� $O[㝾���c����T�r-�A[2��=O�$��cL��zt ���D�<F��U\M찂8�����W���vԠ?�΍ҩ�~�����殳L����K���`4�A.1���ҟ��]>{i�BϚ���<	���;�
BJ��f3��H��)��`��z҂l=�$VP�10#���$Αw���L.Oi5����ۢ���i�Ѭ�]��;>%��KK�"�1�������Ga���-嵕ϸ`1I�"��_iΡm�i�^JpF�q[x�|�?#��x5�X�]T�k��,@5l�Jo�YB�ob.a��wC�����Z���/RR$~w}[NP�=*2�"�10���օ� |�D����#��X��{qz
'��N��W2X�4�! �9��U%�J	G�*(��֌�ƆP8Ł
��Xԁ�n�{⭋�Z��pl{�����$�וG˸7� �B.uX�8�m��l�ҵ̃�T�b���	i/	�~�c�Y��ú��d��KBۋ�e�L:zN݊�K��AF�!�C��s\~���.�7��9>�⵿Nr:���i����{�P��̚��BG���@`�,/�Q��&zյb�t�h� �������h[P��6	�Nۆ���M� ��㿞-��^�ȩ���ƌ�Z�%ڈ�ڮ^n����4��%����[�NN:ײ�M7~���oF:C_-u�����t��L�?�|UEb���P�x.�����)=�L9>X��+�B���&�|1rO�@c;qO��4x����]�r�㩓4�m��H�{�/F����ea>����K�И�#����Hݐnq�0��Ҙ��
���(�Sj���![��|���eI2o�,u�:��:U8�<�UX��k�9M�|QB��i�i�?���҉�<�%�T��Wz��I���US��zv ���?~y�Y�� ���db*FE=��Q6e���ϒ�J�)*��ɮ��70ױI@L��9�q��}7c�ݙ���g��N����h�7S6mV<�&���n���^j	��������/tC��t�KA�1@����$��x��ѣ��ȴRa�}q3T,����E�>��>�K�v���"�f�"=b�8�%���D�@�����7��SQ�c�u�%�`&������w e�4�PK��fh��b�4F���I��?C����F]�� ��.A�cI�Q�͉&7M�Cb4�~�*�fo&^`g��l9��3(t�����w|Md�1{E�}��eo�
�}�c�SK�G��#B,�VB{���{E���! �f����R�'CVF��QrSDd����� �5�ǉ�����@z2u�l����k���6�(c�_.kE���j�q߶� t��,��6X�[6�lo��i�խ�xI�&3T��]�`|��U"�3X*ܮׂ��=F��U�ueG���8fn�����r�\�]L�'	z {s��	~cx�R�n���̟�E���b����n`�g�"1?�m�>e?�A��n�:,z����/�w��vs辝-d�~=�9*���������z� ��`���G
�05�c	���pkpm�r�J@〝�V-�a������+�X@���{Q�Fe�3����b��6�c�7�q�˭�Qz|��XL=�?]�f�7�����)�>ǆ>a�X�1F�:��_�Y�n��L���� :��q�ZC����e-�k��ό�g��a�[�KApWr@�-&�|O��j�����n�x�aƑEPI߽C����4���5+FE_�i	<4g�q��Y�����{���u���ў�D���;���^�x��c7�g���f�z)��$��C�i$�@��@P.f]إ�1C{���LÀrn��`5��C>K��h׮�1 1�A�#�Ȩ�5���~�3W��Rt`�%�RxA�W�@
_l,�����1v��#Ps��2�w�g�I�#S��/�O��8����Hw�ޠIن]g�"-if�}���-%��A�W�EA�_�m��LFZe���|�@�nO�%?��y!6Ն����*�:�^ԑc:��:?��3--��S��Mo_�/�\�����ƼE�ؤ�N��<$��2mod�����������M�����`��ʒ�'0((~�,�+�{W���G� �ǟF�bD!#���̫�N�TH����'�Rd���P�j��A�1�]�*�4���ũ� ��1v�n�'A�(,�iݍ�c�Sn�Q�TNH���OF~U���0��eJ�2� ��O�P40�����tK�д|o�Wo�ɢ��2z��ܤ$qjO��b�����!�I'�}X ���X�hJ�럃co��i���}�u[>��
U�Q�	����L(���AL�I�?�\�͗���?���!o;�������`�vK��A.�#��Ѫ���l���u���!aP��UK�6.Oj��F���~M�=ua|��'�"lwh��-�_
�e#T y��з}�+��I�"�f�LVy�8q��n1����Vp��ٰ�p�K����ah�Y;�M�_l�z���-
�_
�(<��]���XlxVHYEB    6184     f80���@��VK?4q�>��%T�3b��<�uL7d�hI	�k�����*D;�����Ø�j�H���x��~�o��<�����)#`x7cOϡS,"B��P��j��j;�������Vd�Fad�f���U�5F&85�G� �W��=��"'��nwx�Y�A��~E�ډ�lp4���@5P~�;�8>Yh�%��Z��hmKW���Oa�1v�l�!�����CF����w艝��H�}���6x�^�ŏIZ<�2b����rv���y��qs�ĢعNh�@_�
�ڼ�@�5���C��=@W@{�{��A#�c��̦�@秠(W�3�;}n��j4��b��b#hW.��.1�E}>;�|L6>Aӌ.�����hf��K�%<�CƂ���~d�af�2�2�yN�k�
iv��߈h^�k`Ϫ3�3��h�	��=	�<�a2qU<�<����뙸�a�|aj�:��Dp�n"k����*Exɡ��*��w��R�'�q��{Y��
���/���~n,y�)4� �R�2CMn(V�9����	��X��Cߗ�������u|��tx����x�/G��w�'�,/8��&LD|ˑ;eOx���cH>�n� 3*�U��bn�� ����2�Vs	)&)䶡��ͧ��wN�+���`Ʈ�e��C����<oC9V���&���>;��M�ͥ.�:F�7ako�n<{R1�)1M��87��+E�-K�/x�� f��U�I�t.ļ�����^��j]�0h!(s�i;-��>�oE~/x�ZWVB�����]�e�7�Ph5��"�*�}���J�T숳c��ӭ�Īs��>�3(�l�p�"�ƊP��v/*l��2�{�H��0�8=�z��.9�����"�Y�e�2�K��k�K4Tĭ{*������O�^h��%C?��%���WA��g
8�t��Ν���
�%�Wݸ	׬؆�oq��췁AX�L�f#�]+�Z&&k%<���#�N�W�SȾ@�=|&%��ga��!b{*xA���a�u�|�2���U�}/�p�2��ST��8jq���u��bJ�n�n�|���U[1��r��}�x �C�	��x��wwĴ�*�kk��3�D�NyN��_�mx `h��|�
f #�2a�"� ({r;X
<�kó�h��3������z��hh�]�@��π-H�q�<S'��/��8L�*�B�5������r��U�+�a%Ʊ�¼(�V�l��Y��6$��`������J���JYoHG1�M�\	^*3�)�������5��A�i�2�s�.ab�XVo
"V��/��^����O��� �麱�]C�VW�<�T�.�[C�+CJ���|V(�zIR�q�,�l�׊-[x:$rT�U�(,A��[��=͒�-P)��	��\�Ύ����:�j_��ik��^��:@]��'�h���L�>W:�;R �q
ܬ,W<�&5D/ŕ���Ū���0�&/�Km_iQ�>Ьf��*ӨȐ��w�jp7����s���PUw�;S,foG��ֹA��=�`����=��y�6Za��A���&��-�h@00~b0�?U��=@&�� y��1@�M"Qj���h�dH�^?p��gѕ��p�z6}�H*Dc疢h5*G�0�ϲ5n��'j��=z�#~�y�c6�4͌�k�2�d���~Va(��bF&�QS�Y�r>���ȨZe?�?t>�DF����"�_����։� ���6 %�%��nU���*��,�f9��8�9K�hSm
���ծЌ͉9��G�o�|���T|ן>n�l��W�U$�cCS���i5��)�M���%$�w}��qZ7C>7�4�>���??�y�}Q4�� f��s�Gå��L+vˈ��S�-��p����|1	��na_a˕Q"�����؏8h��j�s��%���s�v)�����l��S
G�&�=pk�R���
��L�T������*���p4	O�n�Ǔl��A>G�"�H�`��me*��lA�xCn\>�2ra�eY�J�B=�>fN>�W*�徲�_� �q��?�y���4-j�Tղ����a=�6Ol��P)a|���]���"�pGUC�� W��=��oy��Qku�h��]�X��xG�O �7p�ۉBֆw�aE
.�����p�9fU�9c��T#ne��&�TJ?xŎ%h6�Fc7�ǌ>�hv�Ȃ/�%=��м�n���.R� {�)�#�&q�"� ��>�u��B䟈8Sz���Z�f݅*���lϼ 둤�!���PLŰ��s�D��1Pf*�;6g�P�VhS���_-&��p��(�O9v_�_�('K�C7z����0h�!#Do���E�k�*���Ц-M�l�a`���e?��F���?�m
n�x& �ړ�G�&(��&
�K��xQQQɧ\;���(����2>P��Q�i���'�Ը�N�O�� ��Ȁn#��XY��3�,vM<�j���M=�ؾ)��M��� �̘Ƕ.On}�#[�LL�ew(��*:�9�݂v�z9J���AA�!1-�DZ��\w� 
mYR�ۚςy�u�Ds@m�61���?e�4����%�ʓ��_�p�tMH[lZpV$�Ӽ�=ٹ���M��V'MYR�Wo��K\�U�gT�b�E����w���S�i寮L��d:�*e��;�@��P��� ��==m�ތ���M��b'�uG�W�aȿ=J�=�`�Q��]���4�Pl�w�l:7��C�Ӷ�\���>w"M��K6£]���Н��[�A�Oz�"�bT�|���f��&�R��o`Cb4D~�^�bw:�RiԮ�y��NdE{#�\���<�s-���n4okho���;��2���l�+�0�4�5�����Z��> <zv(u�;�_�f�0L�`�1f`�Ÿg5�g�=x)]O��v��x�;�6^s�������qzl�_���DYB�l�v�Mtr�^�b���4n�X��h���w��o�CP��eL��v)T_Fj��V��g�bJ��0�1�\�h��L�Y'I��8�ܞ/Q�s� (�6�ŵ�/���=�d����C��(�m	9a.�Pf�pa����gX�ި�5�� ��0س��Cd��%��O��I��z���Z�PA�opJ��bd2�=�GlĖ��^�(]�[ /�i�_e�osY*�[CF��˼+m�r�4��dڗJǮ���Y/�}݂��3�7>-ҙ���|�S��p��,���nk���O��S���;Ȱ֩��Uf\/�dq��&=H�4�ʽ�b�/�2�wý �Mp��՝ G����۪�k8T��e�n��a���l���Ǧ���
#)�O�P(O��cRU۝�/�sCt�����P���?k�N������
���
���*�$'����i"L�ȏ��o��A �*�5�+�у�����_�E��"k����(K`.s�[�w8��ċ6&�Ts��+���#{���C�pOHJ�DCә�p��(9�� �}Hߓ,)M ^�Mb�;������É\'�����vfz�p�nl���(�!�9m�%��?��]���Ƶ��t$���XH���
vM����l_��M��4��u�)5^����L������O؟�!nnYP���@@����c��D՚_��7�e��g�'M�2{Qj��	
�!�()�����e��6~r��sk��㢏��+)�r��輠��i(YҪ��Pt#4!�B��
�:�i�d�gʠ�Oh������L�̢{'�Բ�Е贞�~C�x����%W���|���q��M�m�w+�IxMW@��Û�5z���=�y!����ȼ^Y7b[gp��ϕ��q�'���.r����1�> F�t���R���KCz_����7���u�