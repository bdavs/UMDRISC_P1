XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Fi渳1
�k�+"̆����o2�^$6��kQpO�ݔ�j��
�Q��u���`����ޙ&|i$���U�_�scݧ_e�+2�#)��ZW3�A&�x�ʎXnbҾ��\�����8̚��
�ghT(N�$z�(�0��E�,!A��3�{Ϯό��Ju0Qv#��QٲT����>O6��1��2�-6`�h�G�kNۈ�9=!�;�4@dXh.�+	�0�;�:������ō��#�9��H�(�S����;2�w��٣�����G�#�#n�5�`2�o�'��A&TEZu�cbC�gk�žY't:�"4DV�yV��j��j�K���毨�˲U��%�GeR�e� �P��k�jZZ�0����$�_�qG���l�@�nP���1�[8��dS�>��5��Av*���1�|��$3}I�-��f�l��M�=E��J����#�����p6a�E��z�\�.�/|��v�k`B'}#��F���$��F�.�b;��v�N��v��5�_��3��Ou)�",���x�]���P�������-ʰ�͂�ㄫr<��� 戓3ZdI�*��N�I��ǯ�V&����cgR�3m�P:z�^u�@�6⠋��6��e�3*za��*�/�[��2�S)�,dx�;�At�zl-\�/�D7g.��c�O�.�Rܓ�zG�1�"�!�n򆠙���3>IJ��� ��}\��.���`��"�,-�{�~���~��s���.#��_Q�SeI켥�,�ğO�N<
�p6��#DXlxVHYEB    b631    1a00��!�!I��J���/r�г��Y.�T���-m٨x��Tk[�{Z���	LAEt���T؃��r�o^o�C6�#��~1b�Vs�X`�AE�Ӣ�;Zis��?þ@~�2Ԩ��9����~J��F�S_X�,
��{3�k�~Rǻ,ғ^��9CTD9C4Sdа��R)T��|�qV25�eR��4���!��瀅�`�$���'�e��V��Χbr�3���<`�a[�_x�]S���HGx�h�Qc�~s�rg�|M���gh]���+cM�r��]������ñ�jְ�q�R���5��a��ϡy�ċ>ߡ@��~M�tu�V<2��C&�+�,<c:NgtHT��4�k����C���:�iӟ�D�7���a��:z�b$��V+�fh~,>;z��*�� ��Wm�s)R����0C��/ܺ�n�z��^�=J����>/�t�7�/�0��~P-�u;�L;����Bؐ���@@�[Hdr�E��	�e(�s4�D�Y�՛t�ro�1>mΣ�����I����G+)lсW��hi�q%�J民��w����ϵW��hw��e �j�˝�kY�G�n~���;ܓ�.�%n����rj;C�����c|f��_����ia|�a$t�ޞ��iy�������$�#�N.�
mι��G&׫hU1�F�)�g(p>]������v��o+��;��'�۴��o D���F�hz��7v�>�~��40TV�z�+�V�y%S5X[RVbe�LP ��i���M����[� ��P��-Wr��{F��O�b.:���3Ѽֽ��Վ�`��O��>�we�?!\)IQ�%%�~������$F�.��򅊝�bp�:R���p��y�@�rs��dS
�hf���ss�\���YK�
����(Q�V�C�[s��Nw�"��Hy����֭!ب�6C,ԑ����ϊ	L����~Q��i��ls-��}�+��ߍx���Vi[�EY�?���\e [#���MgN���&�̝qOT.��6mD�O#z&�en����H<�b([�1q	�^�-I$_<s�1J�^Fh�V� ����`�&[���3�z���NN;�V\h�oI�	dg�������	������x��c~̺���g�Ѡ��;]!�l^�0�A|��?TH�S�}_�A�I.p� �_���~�]��4��RQdKWRwm
$�Ô���Um(�H��C�tCf��q)M���NhpޔI_\35:}�\~�BjAڱ�������C�m�4� ȪG��t�Q�T��aO�5^Ur�_0*u���o��H'7�C����TG���cjRp:���0^f�.'"�2C�6�A�J!
{�^C,��l�˾Ɩ�F�� ��1�4�K��5�w�z���2)T"�N��*�N��$�+
@TW'�ƞ��B<�D��N.����QE{�a��т�£%��6�3u�E���c��\[��M١j�>�\����'V"K]5��S�&���!�c��������hu�!~Cݞdq�͖�_���Y���4y���kb\"�mw7^02�','��jsX��̺\���։.r����JB�ǔ���L��p��]MDp+�O�@�,U�QS^qx�nVj�!3�̔#Ұ,Ӹ�ܸ�ʵ�\�S�DK�RShњ�YX�r7�H?����gzk�rG)`YM��Øw!+�'�^�d�ŉr:}�>��.h������<M?e���)as�[nٱ �3ZwV��{_9Bv�(�"F2�����
]LrR��g85�T�ns\�%�qS~h-�8b��ݲ�wx�C�kY�'����^}�(�!���U�F}� +����6դۚ����ѡ��G`b��=��s���h�c�{*��%.y��F�I�T���=V��{)��q�{]��j��lY�j��1��
0��7�ق4¾u�*^�vw���ڻwM��U���
d�.�l��8���(��1����hcl֐g��@hCC��"p.�K�¡���XIŻ��"����A���-�߷+��7���I�K�!�V��D�c�����Y�#����{�܅"��ӗQ���b���x��x��(�c�q1�X⪻|�[�6�."�ə�w�2�ky�p��1���d`�;���� 9S���|� W6�Rs���	Mѝuo�E����^|�6v�
._&�V>1fo�Aߕ���""KC���0�0��3�;��?M��������e���~��?i�
����Ⱥs�Ccz5���{�ٞ~��سx;��	�,��1tq?��eD�������e����]�!.z�	ǋ�3HF%q:]J�YSj��'Y�[�w�|��i1��J�ӻ����o�2>���6,��
06tQ�}��SpF�p<*�~�_��V��&?��I���t�8e�S���
!.�j%���C8�IB+�9��t{`���d�oW�eJ�+���&zV��!V]5���ܰ؟Ji�p��o�m?�v�Pp잘kv��t�s���A��Fx�e�e0�3�q�� 2+��� )ΰX\�_s�3p�ycz��&�J,������\\W��G�%z A1��8m�P�g�_�����K�������'�R�^�|VҤ�/�GM�i�\~W���7|�p�/jr�Nr�����,!���;��l�5� �ȣo)J܁����C�|է���E��)m�)��6Oׯ��V�M���8*�L��h]W�΢Cq[�x��������E��8����k�̫K &�.��_<M/��k��x� �}��+a�]� � O����*&5j�_5q��w���O�i>�����!
TF��PW��E)�	 yŰlD5R�$�h�>y9b��������^*�8Ӡ4�h@�no[�!�K���,꼩�5RL���
�C<?zJk]�n�u���Gb^𤋮�|��]'sϨ�5�!��8�����i���x�*I`n�mى#��=��:�확�ف���t�vl�c�J3f�+`��߇(P}D��D�'�8��5� �q#�� @��Xb ,����@Ϡ���9�KIu�zP�����h�ze��*��3��Z���@�}=����	@����aX`�sJ�{�jN�1&ؙ;�D<n�+Um�/��8R�f�3�B��h�?��/Ť�0<&�^|�z��C~~XAWY��*�e�"�O� U-y�}�{�����'�&ҟ��C+��d��~�B?<�u=ߜE�~�?��I�B!ւ5Z��Δ#?�h� �dK����e��*��ח���U1�����	���M��A��������I址��0�0 �����=��!(�5�g���?�"�ŉ	�Գ�����u��T >��
��ZOك��@��!�p��n�l���_���s	�z���$��*��Â�/����|��J���>�o�����M���ʏ�=������NL�4�[�p��IS<�ݻN�k�;.�g��j0R.\�����ΐB���n�i�H�#����v������5��L������-d�	���]Ko��{�K�޿��$ls����O^4�ha�W�v~�ieG>��#i[X�n\�*�m����ph�������X��M.	^��7����zkiZ9լ��c�@ryam��h4J_�XtRx��������(��Z�啕�k�7����n|�
�r��0����Q��<ц
��[
��J��kH�Kb-����Q�]������� ���nB��^��j��Ee`����J��<�KE����*�񻶡��g�_oZt�c$�OLW�"Zxm�,�7+�+s0؆��K�mmF���r���i�5t�#���b�Fױ�$�#�]KNg����V����ZM���r����,Aѵ�~�:.��6�i�'��d����:�jw�"�i�S��3�3[�m3B��\Vc��u+��.�ȩ��ؘu#:���;ds�fH󸰏��a
|���fn�Nc��n�ƫV�m�_��̠���M�}���1`��s�Y���ΧΠM�Q/�[�a��C��p�p+��#c��.�1\W�\�XL�$01�ۨ�[_�ݷ��c���v�wNI L�^��ϛ:���u뾟�P�dAm��e��Db���B��S���>ӛz�s��L���I���M珖��94<-��tsۦ�rh�M)Y������gPZI��mރ���9�6�p�`XoW������8COߦ�%g�bSF"l]�nN�G�ݠ~>�M�j�"�Wa4�(�L�w��e��ʒ �٩15�4��X=H����e��,;4{��+���`D?��4Ȱ8�#P�,����T��k��M�����l�j�IN���"W�ö�I�9�o�	��HLK+��ES5{�D ��P �|A)���u���C/8�-�dZ�Y����ꔊa���OU��K�v9_P1�K�Uc��#Z
�~�wy>�S,�ճͦ����:(��"`b���`Y�t5s-ru�0���-Z����h�>��%�5 j�ZA*���֘�^���=��B�Bp�29'�����;s��A�e��;%��N*]�h��� ���� ��7Jm�v��Wh��̘�x�ҩIDu���\��X#��!;�6θ�h
u4�b�[ֹ���d�ۥ���(Ì�z��-}���)�F�J��BEh�[Ʉ�����򶼂JO#�����v�klE����d�n��Œ<�ޔ���b':D+��,By`�h�U2m���_Cƿ���N���h�v9� a%�9Iq�QS�S���^��Z���<'=����m_�̀�̳�8��⨌�&� /BC0��OD�߰�r?��J�i6 9c�g�`$�8}<��������;|�sa(��M��������dW��P 1Y(W2U3%��^'�0;��E7���d��)�C�p�9"o�i�������n��}d�Mf!�?�>���,ל�G�P�������V����pKHNg�����rQ���٧X=13�b�W��X�_y�؅7˓��-��O�3�R0�؋`3�[V���s��eƐ2Ke	\�s ���Z������,���M~�`t�f���<N��|��G�O�����.c��+�8�o^n�ׂ[ݼf@��e!��o7]%-h-��5�܏����@�!��g�K,_�RuL���>�=k�o��alyd�ݭ��hY�?ޠ�O�³�u�}��̝&�z�*��/�OPm��hP�=��i�C����%���{�s=���3#6�u� k��e����u4y��������ۿ�Pub�� ��S��A}h� ���Fa���#b($,>�g�t�������V�j��T�G\���7�h%$H��*x*�t�H��%N6;9�������@��X��
�?���p71?�ܾ�L� x+=�F��̒{1��RyiG q��Vֹ:ı1��B�	Мnߗ`�>���\�'F��� Pz�&�U�� 5ii�N@d�d �<�Vܩ)��;�I���{g�l��2w�����X(ɮ�<��RE����������"�i����*�>�!K߷U�X
����z�ӌ�Bƻ�G�\f�1��3�ɷ=����'�۬�˜;߹�Y�{�f�/ַ�tKTŷ�ef�f&t=�vĮAolF�����'3�A�3&�e��!i�A���0��ENg�uf��.XR�6Ij��z������E��SpF,�I�h�+m�}�}��H�<�ZhbS�zy�i��J�B��4%kn���̢���X�*AN�K�u#���򘔬Q��t�aS����J�)(E�)���DC��ɢ��F�7���� �+8?������7���Rh��Ā`I� ��Ri%_T�:
�F�ژaF�_�i�0eCy����ٍ���X1��#P���	_�^Gi/t�t�	`����e�`���˯�$w6�,/y���s����3qI
�����2u�Y��;��1��_�q�c�х2G��[�)ڇ������@]`��̜�)i�3,LOR�(l����Dv鄎�ڷ��o��hѧú���6�s�SC��k�k�p���Q�sz�:hAn���^[Q�'��]�T+ť-��ҥ)}Ě�yn�l�i0��VP/,m�,��L>#���U�a���+�����D˘]�h���[����#[�{*P�`���>J�u�r�S�:wl˩S�*����q[������_՜��b u��B �>T5��irFT./�t����d5��6�Ô4q��T�I���m�f�Ǣ����"�p?J'2�����J�i%"��^r%����gK��F�Ll=��(�:�]�y�юϔ�1������h��^���{8�i�����8�=32�(�I��x�I���^��|'Gu�)DyqA@�6��
�䝈&ٳ`�9yA �,о��+�qٵ��Zƞ?']�}C�#�5�))WB�4_Ui[�*�gro׈�;�����6Y0�$��k�<�˥��. �un&�B��	����&�ZV��2h&�������gd����EOW>��`:��K�񖌇