XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������O{[�?�=��8�갩ϮyW8SX�$�\(,���k�*��DӺ��ij�����}Ne��I���:��ΆK���3����B��̧Z�},i��U�ce�L7�V�$V�Fq.��:r�
#S�5J-�,ϖ���~tx/�&�Y�H8�DX��;TӞ���-�<\*�j���i���ȑt(�}�jk���r��231xM,���*xi�1����D���#�ᰧ����RS�F[G	��9�)j�Ӂ�xC,8�ښ��<=C�:T�Iі|�D��P��,;���LkL:�r"�#?z�y��t�X���WbO���Շ�k[|�E�����/���c�;'_�o���U9v��(����b�G��)��1�7���W������V0��&Ď�E�Ӧ'2�,ZC�A6���YE���a��A�[>�5 3p5%/�����zI��.� \ȱ���0���)災9ݷ���+;�(.��/Vm|��{j�X�D�S,�u_��T��� �t��x��gB�����i������3�Q3�;�"�ah'�����b7Mr@P�^l ��0�o���A{D�?j�Pǁ%�
�m�.�ذ�U�3L'[!���<׹e�������爊_N��"��}5(qF)x�{&���ٴ/�F�`h-7�7>���4�����uj?��'(z8"'!��E��'�(�zX�Ü	f�8}���ťЅ�0��.�Ѻ"�5��}E;��hT'_�'��Rkӧ�%�ׁ�w�<q7�%֛�ōXlxVHYEB    fa00    2020X�CK�D'(w��U2 �6!Z�@i������>ޤ O?*���_)�(^d�˱1S�3>h���y�(��n�o���0�~�Ĺ�ג�.���������R:�l��ĪSL&f�e�c�����«#�S4	 N�2���.�\�%vH'����	!�1s�& 5(����:���)TO��H'ķ�+؅�T����{���u�BK��ªg0�{��`�ARBr�!n&�ej�HEr)�YԂ�ň�d�<��@o��H��f~ �F�A��h��~�� �]����z��Mpt�Í����>�k^���=���ПT*jЫ�o��kl���h��������j�}�bCr�h�a����N�Ɠ�φ��q����̠E��;J����%�?��-�w�y؏DIAv#|Q�u1��\�p�A�_|#��j�`�{O4��Hɸ|��:�<��8�:k��ա:�OXo���s`@G���X}�}�9����N�~����g�� k=�oK{�A�����K�V��|�:��.�9:��� �k[�?Ր��ڈ���zb_��Z�"��-Ӳ�XQ�E̾ �������!*Ȧ/�xE��]���\��mW��:�i �}�ʠ��Q=c�%e�ߧ�6LaWh7���t�@�u�Uy-�����!fvW��c��}�@U�;��ɜ�5����Fͥ�x�4��>�'o�@� ��2�"��4�MP�<	�JH`T�G��Gɵ��4�38
�pgj��ff�\|]�Y��ǠHcG�������jS؆)���=x)��O��lݮ<I�	�^�0��gݛ�!�+�a��3�<R����'\��iE�ꮁ+��}.`�} g+�Y�(����S|�S���fB� `]�~��w�ӣ?I~ÚG��W �β~v9v��-|�=e1&QIN�Ox�r��}��H�=�,��m��jZs�jRVN���W�H�t-D�j�����5���/�)5��K>�?��ȁ�W�FaϤ��x��@�m�J� ��Wv��Y��jy�%����'�lIl�W�!��H��Ѫ�/��me�������ߗ�&�àkȻ� @4٘k`7ɐ�s���wJp[F���۸�3Gl]����	Zv��1,����y���)�	0���`�u(>�j:N������'t(�.�Cw-O�p8�7��{օڍ�"�Q�aZ@��N��7�Iy\���(ݕ�z!U�۫�l�3�ݸ�1WrCI�b��'z���ƌ���܂���������x�5*r�׫"T�jW��2HYCU.~�Zm�)L�v��U�ؙ�S}���LY�,��x�:����1�m�n$ 
�������w=��s�U��)�
GH���5��j�#?���-�ֲ�V�p�n��8��{���M���:*��]�uf�G#�9�g�E���t|�r{T;���}���l89^e�
a "YQ(�F2���౦�wD��N����(eI�L�����8^�좂�=�p�9׊oH��ү�bw"�BCD&�H�*�f�X��3Z]���vq�5�w=:8��/m�%��XZ���{��^XB��V���ėO���>�tD2;��F��=�n���D��9ap�J���-�B`��{9��h �����:��M4�s*��g�$��5���!���l����J�T�����f��&�s��_���ړ]�-���y�zJK�"�ӿ�_�=�R�?[��D�=�{����Y�W��l�Ҡt�����0�?nHĐ̫ZBc��I�Up���N�!�o[-��|��#��!�]����=�)U6U�.�O����]�^���p!���Ћ?E���0��N��]\����T!�5p�Z
t^4�|� �RV%*�k��}��V��N�G&��de�/�q�+w����E�ݰ��_ǁ_ ����@�
+�@H�9��@�I�m������h�����G�
�k�e�d�\��cu��1��b�mS�W�/�Q�Y���)���+�BP�r����1���{a�^
���{���z��k%ޤK�@aY�}#�;[Z7{��ف�Z�v�X3,��SNbad:҅z�X��m�~����>���i���<ԩVl��p���������>a��k�i��d}[ 3� ��Z�j�x���c�3ŉ�:�agZzn������E\��6Yu��)!v ��m������|�ҖF2��	J ���u��QNN	��&e�2Іr?�&�.?ſX8xF'�LN'�U��z�B6Ғ��Vhj���0�v�u��g/�^]�
���p�ĦF
�ZG�U��ο1��"��K�hjJ~'������CKUܫ���2f@��R�Ν[����ɻ�]JG��
>��2�*c{���f���]��������`����*xn{Ҙ&�Z0+��1rC8w�R��=RT�bl�y�Wz��&[�;\D(��k�0�=��a+"I/>V��� |�Vj�*d�$[|+*���ʢ@�R��3��b��-���
�ۉ�٢�;�h�6,�EY~���|%^]I�&�Z�8�Y��Oa{�&P� 鹎�Wpn�OQ�����7Q ۭb
��ȐS\}ѐPvJ�%����¡�����4AШ�' ���@����>|��k��x�R-C���-�Gj��P��Q�`��f��。��Hv�RI�V<�"�A�}=d�F�~!�!<9��K�Le%�"�E�Z��=4tze�K��i�'���9ywXG:l���j�4���{��	w���c�I\���0�_^���o��_�>�q��j����'Z�H�U��[�F�B�䗒/��3n�ݟM��Y{��)��A\&]*}�.q���䏵NgN�r�OF��=�B�4�lq�	���{��7�hZu��2!��]��0���f���P�x�Ak%���N�8�x���Y�� ?N�3	T��I�S�v��.P����Z�:c�k*��wϺ�׾�,���<F1z�jB��o{ҹ~��?�IK�ķo�c����J�:!�q�	��$E�{(C�	oV��?�S��E3��-�&Xsw�߿[�pO�p�v��8n*��Ht��k>�/i4���*��61����;�x�>�����9�(0>�ƔѷF5|��Z�V�8��2�*�����)�)b/�1���9�Wy?����"!\��s�c	7S��z5�b�<B��0\(��;�M��.(c_D��$}6c� �'��`2�>O��M�=M�C�WF�lRR�� �y�tP�2�Rq�Wb��XS��;y���ɴ�^ +7����l{�?M�x���ʠ�O+
��f��5�=�qk��4ڶ�O�1���� �MP|l▵���	��*P���r	�#l^�"T6vU��X�u>�Q|ߧ��%�%�,�P�a.�+ۡfzj4���5��^��]��G��e��g�A2׈V���ǻ�`m�K��(�
�vZ������{�K��}��O&?q3���9P���C��p���F=ئg�;��-�ė��b�-�a��:��?|s�#���Z$@[Go;��Y�t+VZ�c
}��~y�`C�F��+|U@?:����cp��.�[���?�=A tLƫ�W�X��([/pa�➳g{s1&3 ��@X3��i�%,�˯�bU��jt�6�Re;�mX$Û�4�?/~bZz��`hHGe��v:�ą*Y�cy��zNt㨩^��@Ǉ����'R4��j���@z����ڳ�!�T����)�O�ہ4�Vm����l�w����<�,�J��J0y(����_��F�7z��>����V,r������Ɍ,eěU�c(甤tU1)����Hb��(ޏ������ݣ&
B�&�e����/n�c[�w�>Hm�4���R�K��H^���1P3ٟ�|V�/����c�!"���T[l�?!ç�4�Ze\_#�������l����J�_KǢ�4m�#򠽿H�:�ƭ8E��j��*���~	�Eh���0�����ՠ-��5�!ŕ��+$���!|F���x���W{��Z��� `rn���wm76���$�*&(��l�V�&�Z�A���l;��d=ER��_R�e�8�Y4B���'B r=7��� ��[žÀ.Z9
[�8�+3R[�4'	<��/R�-����� i���!��1l
�wgXpP���fܟO���}��&esp�
�v9X�qs�<���,�X7�H���n|�Ł-��'��"�{�8��Y��f��.oe[�_�u�|O���������|1�,�t�z���9ݾ�L�t�r%%x��"-,c��|8��;@���V\qɕ��dT.ÌyUNWٰz�ŗ,!�*	 Y�`�:$#��C"�U�6����'�� <aeZ�gF��ς�g��)6/�/\w2$V���aCH-�@�k�g�����w�f�{#�[4T��>�m-�~$��c��̑c��l� ǖq���դ&:���<5�w���4*c�A��ڞl��Bi$���DA#���V	�c��Amo�m��ݕ�c�ܗ�����d�w�5��F�>�9�n�E���R�E	�����ᇧ@%�PrK}|QUI�v%s��EB��J=�F��:)���L�㇎l��T���~��hpz��
�}~���et�;�ٳ�Z6�b��&���Q`�(�L�.p��"s�%���7aG\��z�@{Z�@��Ko���J�hu��E�!C��Z 4��݂�v�6��Gx!�K�I^#����8OkT���C��vፍ{�������(�1���r�\�0-`�"9/r���`�̒��!�,������������Ld�����?�	AV�,�ŭ\ir�JD�Ѐ�o���M]�5+|
�k�X��j@�7ĈS�3̗`���gg��Yr�����Hy��L��7�)R�ș[���81[�$��]T��>���;�cN����B5���ى*�V�,ޔ-���N- �`-A_�@���FD�24���������*i�mr�M*_�����?ì����Y��t�.��A���x�d��φ�b ��#k�v�����l� bU$��Z�����/�F{�!�;����榸��@L��Т�/��>�s�� l��EUgB<׃BY�Ey�h9<X�;�v r�����$kҵ�+X���k0K\~UBa��8�p�C,���ߋ����@��l��ǻC5��n��-s��[>�7�.��O�9����ʏ�"�u�/��k��}v�#��/_���v�� 捜�)��,"�%d?�>8���o�g`����6��j(�܈h�b5�o�`�Yz�=w�@W�ڝ�b��D��-	���l��2�_�� ��nK�����Gw$*��KzA���$��i)�"�r��؟�C�a4��)�l��<�2֔�=��W�\[
#>V(��\t�&�+!�iL�@r�6��Ht<�W.�a	>��U�"��w�k �ɾt�g�zwV=P������ 7�O�;�Y��nT����'RDV_3�'ˉ���%�-�{P������r|�ق��K-s����)�utkĕ�0ڑsٗ�HQ�M|��"D��*�_8���D���ED�J������t���I��q'6;R�'!`�B"�����;㤻�2�e���u�'�h�����nF���"�I�NAV��+C� �]�o�#*Oi MP���ķY�a:	q�t{�������1��oWB�M�`����s�)�nQw"�[<��Yu���uC��ɫf��FC��?��J�za{v�����EhrΰZU��&�0MR�Ȕ�1?e@,G,t:�����XЂ⺩����G%�EuWӉ�ϰ�~��,k�A���>�	<p����9�b�V�%j��}���sn�NLc= wF6x�r����ߕ�-΀Q�)~D�Xr�Y%����� k�t����� B8�&��&
&�{��p3�j��YZ��͎H��D�#A�V6Gt�q�Oa���4��Sv�6u��Q��ƈ��F,��T��$%��v�n����u� �ب��/�Y�މ�꾘e��i����eJ��+CJw��*�:�U�W��΋d��_�f臟�d�'x!�\FV}@�+V�Dx�|#��,�|a��4����~��0{$���=�:��Ǚ��߿:�QZ^[j)[�8B�4ܑf5hm$s��F���q��^�)�/ZXI}�o�J�&�?$!ˬ.I�I��1w��pD��"ZSn�tN�;���:�g�b�3y&��|�d�%�N{�� ��׸�v�W&x�kƟ�z�B���iQG��� m�$�,D%N��sy�ˡ~Ù�S�`������R�H���-G�)�����dh�w�}{s��9��.kX�&r5�]N�Y����kA������C:��(:LY��{����9f ��%k�0�/��̃| z����C�x	�����MLZ|�C$�p�p�q_LQ��z[�Y>ST�e)�?��삛R�&����$D�e�
��s���<��U����VG\�ֽ��LB5��\e[Ϙ.�C`��P�?���h�O��P%�;���1��@؃��U��f�sS�D��J}��.X�>�^�6蜡	��KeN{�>��+����L
�\n���Y��X�� 5z`^ ��nM �e���"�ᇋ�&H�Q��L����]�C��Bw<��K�1P�B���ʃ�AU�J�嗗�fG^1�"sA��9h�J95_fbM�{�l��)�hVZ���ff]a�΄F��	�6.3=U��\�%WK;
m�b4v���%�e9tmtZ��O���}w�E�`���*b����Cdg?�Fs�:��o:���6͚��ܼ��_j0U ���
��! ��
�?�'w��	g�K[t^e��OA�.��>(}"��Kh��T�Y�g�2�$�W��rK�@�xKmn^'60,�E�V��Z<3M�p=[�wx���Xv�? �hS!�� XK,QP	L,j����J�cz&.ԋ>�\�5.?�Uy	 !|��(�T�O������(��oc���zm[�'��h�kݪ��H��t�T�H��]|��)|8 �$Jt�#X���偐X���^�NN
��&Fz��\��v�|�)�pt�k/������1��Q�}�>�t��\,t*�d:����>@��*��\S߾����]�Ğ�Nt��C��h���;-�6@h�U�Pz��hL���_j&���c�WC��6�.���u��/6.FǏiv>��]�r.�%O3�C�_|Q��ք���	}��TF���Q+a�A���e��C���#{C����J)N�G:!r�-�^#�e�b�߸�q�aT�}�^oJ��?�>,���*��C+�";Ԧ��)d���Au�
:���á�B�͡v�r���,Vz(?~�`���.�`^9p�?G'Aۃvƅ��Ĭz��g�8����s��D�?@�Jo`dvs"��� �nb�ҳN�W}��O_{������UsZi�Q���c ~�ǒR�_���z�9������Q��*���<B�j3^�n�ɢ�\G�����l���\p��VXj�;�'��-!����~pRt�5�3���%����p�.XX�Ƨ�(Y~�ޏ������*�q�J��Q�{!�Ak�&�^/��(*�̧K�,$˟��vo}r�oڞ$��j��ypb~�Պb���oUQK"5��x���'�����T�,�̤-��k;<K=�:�oF-�>u�J�QK5�ŵ��;a@�0��=ю�K�}� 3�7��gÓ�H�M�,���ɫj6�XK��	��N�k�A�]i�����<��v�K��k�$z�z3]6��e	LX���'q|	�m�Nڛ�66~Λ��_��l�� )������L�,dt4ph'L�+Co+��D�7(��	K<�.H}\C:;E�@�!��O[�bH��&��C�����~�.R�ѫ�.�S��xH���m�aSB3*O%�eS��O���v�:�Yp�2��W$]A>�œk��$�I2̼w���9�Ol=�%�Dd˸[Z��D	���� �%H|�T*���>�*�zA�Tj�ݚ� �6[����P���o�x��=���	���s{ː@��wa=.�� #@{z'�����]B["n�Q�_@2�u�q�SJV���XlxVHYEB    cb82    12b0�'��Mk�.���/.�.��W�Lߍ�:��=sm� +�ΖmC��_��v�ɷ�q{Ô��CQٺpj��C�J+����}&Զgy�e�Ά .ъ�Ex?�u*�Q�Z��齷晑��5M\��:�5�UR2����O�Y��^���]�B����p.t �;�Qn�e��r r�ey�)�=m$�)o��1�����������u�����`�s�ғ�n��OF)�ߔ��K��t�Fv�^������ax}��U4,��ә%[m���e����'�E��q�R�_Yx��J�b%�'��4D�]�g��5_z��C����f�$��;{�Hg����1���,��d/���U��? �	�ԩ�J�%��a<F�P"�<�p�x�*���.�[8�I�F[�~2��P%�bR�;���X�q�u_�5���'�ړ�Ứ$	���#�4��bLX���s��M�5�a��@yb]���g�,)~��-I���zS�բ��X>�I���:�����Wjt/ Շzv��Qv|?�4�o�N��]�)����.���p��y�����S��h�Hp�l���&{��*�����}���
o��L�dU���/ʽ����J��t�ʾ?HB��(UD��� F+ź��׶��XU+��a��C�P�޻}��h|�]v�H%�n��^��'�<�yɥ��d�ÚÇY��͍�+1K�	@YuK�a	�6���%��k+
��Eh�HHy����Xw��H��2��^��v��=З7��X��0����Ō���JFHX7i?��=���
¤��T��ր[��i�g�\cJ��MRӀP%b��5y��tU���]��8[�q�͍S���9ʭ~x��Mݵ�`Q11��
��*>���\�f;0���] ����1����)u�j�S0ڤ�-��O����.P �ڗT䉖2����M��b$t�rŞ���چ��fy��]TB'�}د͠�Ģ����o))(F�rT��\��g��i �_��k7� �@7��U�'/��9m����˗��z���Ѯ�`��A�-{�"����
��W�;�S���ogH�#�Ziȩ(�ZY��c�%��Ae�RɆ����ĐTι�4���\0�lu0h�ٔ��,�1�čxw��{��jH����v$vm9ɚ$���m�ZR%��U0L�n-=[�	R�ة���е���})�W��^³v�*N1��[&["1�����B�q����R���]��e��|#���ҧ��F}X3-"efJ1�P:AU�V����q�$+�c��<y̝m�>�Yi���`S��o[�q���PY9�����^Y|���Cg�ZP(/��y�^��W��H�bE�B�R;tK�n����O���Ծ����×W� �u���Tf�yE��T^���M�PV��ٶ�U $���6D���l�nH?TX�[��p�ğ8\2���H�36h!'�D���|r�OqeY��]R��y�y-����	6x&	���ʡ�R�"�=�O�X^qd����$=a3�Jt��ͨ���Y[���>��o��>O��!B�љ�v�{,Nly�g�O��T����/���d� ��,c�V��9!��e�L�;П m��=ݳ����N����ΓFk�ro�CA[w�e�=�C��	�um�w�sto1��'c��e��c$.�Q)ɉU�@��,�-;H	�R�A�u�-=�����ޥ��*�/�҉��4"Xf�s��X:�[vӬ-Ͱ`�.ϕ��e�y�\�P\��|@��{�cp#�u��B(Ǖ��+iƗp;_�Ie@U??'�Q�PjUE��6��\
�M*���Ts[$:���m�N`��X*iۢ`я���f)y���!e�־�4q�~N'&������C��J"='N�u��wK�`uY�{��Z�~�
&���:Yt�l�����7����9*Чn,�e��vW.���i��ξy�\^���2p�<�]��Z�:_{N2@9�_{cM�O��%��zʪf�{��͎�y��n�?�'�gpZ�;���	/G�b
��D�c�k��*��̕Y>��A
עh<�㈓��QVH�B�
JK�lU�#V�T�a�ߑ�ASzpKV���^��Jh�Z��]2I��h)�Jr�]��g?22̼��`�s�5����`
fq�*��k���@k�;+���e���`�2��څMTW���=�gp���;(�5-+��*28����9�����6�]1}��Q����RR���A��4�oߨ�j9���sK5ѻ��ЛH(m��Pm�{�a�WP�wqJ����v��_�-x���e?Tv��e;�`��guC�
�pt��S б|��Z��K�U��"�7�DS���]���%$�!$�+j��?`�ҫ䪵���ʠ�	�F��_�������r��}���g�Sa�bx���{jn�~�����zK3�[�,Q#��b��1`�g�"g�� � 8�}�؎#�Rk���\��O=;lc�3�]�M<��ػ���5��0����7;�U��,�Y��\��n� ���z�s ۸�Q07�v��4�T�Np�n��J���y�10(�Br�L�@[(�F:W�^���/�?�YI3g�����g���m���6t��Kp��DPg�<O� v���J�q�g��-]0JA���}���eT�C��-JĈJ]�<-{'[�ɨ�eC��T��&F-72��~k�dz�!j�~���76�2g��&�,>�k#��~����9r�G�:�T,�xI�RvB��;�友�uRd��4����~������o�޶�mz�W�Hx���
�i%3�4���a�����EI���������ƒ��Mo8]����{����F���i�o[7j`�z"�>���i���$�V Ψ]�)/����vs�+7�����M�kt��f���>c�ia�_:|�~����?���sb,��{f����t?��t���'��߶r~���Z��i�<w����y篆L�`#w��jw�>ƃ�=���V� ��xȑ���*Us)t˺��1�s���ZK�wPM�����Ո�H�7[&zQK�v܎�Wm���O��C�"�p�0���eOJK�:]�C�->��?�Ū �Y���II�;�!����8�+&ښ�'=����l��B��$��[����0�{��q�'d�Իc��b3B� ��3ɡ|�w��ae���3��>Q����X���ǫ�#J�Geh�}��$�j�el��4ɀ���@*�5-�`>�7���j�+�∸��͂!���BYײ2�i'g�.)� %��,T�Y`)*s	�~��^�3t}�{�"ޓ�>��������#v�sQ��;���qG0���$!W�ﮥ& �L�S�k��ZG���Øx?ER���/܂%� �u�2�
�)�H:蕜X�C������������ی�e��Cg�-���7�G��R�Vֈ�=w{�2�~r�\�p�u�)�V��a"��c�����|�R���!�������ţ�_�6QATI˦�p��]��3nBXߨ.
8�%\X�+)��N5�[n�Vg��U�\�O3"el���0`��X�|�)ܳݕ[q��<�m?n�e�����ubI�}b*	t2=.d<j��TK\x"���L��1l�;zȐ�ʆ$��c���������`K�>��o�\��b5� �<��0zn��4.�{���r�F)S7Ut�=*'+���g����&��M�8���d�CĨ)� 5	bz�_"���â^h�b�(�W.�	�`��uc^Ii�����mD�l�:��V��=��5=�``ʣ,wA�ʳ{�u��s�e��
v� �K�����|)�$�/1�Tz��E�q	���=�����7�>B��&KF�=a��1w�E�(�ْ��1�ڪKtq�;�U��l�~x�"x,��z�y�6]ٸ�!��U3Dfe%*p���Q��I(,m�[0*H�/(+�W-1�v�'f3��\ƹ��8�қk6��/�'��[ɶ�
H=�h^�<�v]7tK� �B�:�J�Z��Z�A�`���j�i��e���}���uy5R�@ɋ�Y��-)�;�&����8��z@.�1z���c�-���E}��0[�²�uG���oc�@���[/��V_U����NI����_��,ϼa �?#q�gu��"6ة��i:��I7p'��/�9�I����o4ծ!�� ��e��W`ufM�+�"�f��`��o�oNX���R���T���׭e;�1q�f�X�k��<>�v���E5|14'��u����)��s��W�$�+�t��m��b���i_y.��k}[���_�H�k=c2,����=�`������r��s��tMr�c�
�m�S�]:�?����k+E�]@ f*��	��#���v[�{��[��,�C�3"�����ՊDġ��G����H]C9����?F��'�����Z��Z�� QrZ�Q5�n�$����ejQ<��u4X�x��7������<�Tp��xi��e��)-�oY�����uRV]*Atߛ��3B�R�i!3`4�2��S��h�ھ�d;��z��e�.T��������"�a�ZQyC�ᓠkZVa֎��%)v�<"�q%$^�_Һ�%ܠ���X��(�D�������ڥ��F���[1����bm