XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���H���A�%l�zм�n$�?��a׆-�ap�����S�0�%������S�+O@#�![����4N��*������t��؆L���MM��ۉ�>UP��Ko3���KN$K���?��R��w#2��-"1�(��0��U>�O�^��u>�s�,>� X�ꂫ��{�)	+M�N�H��4xS�LB�����P}Nݥ�0Ne��>�ܮ)Fq�J
!��;:��f5�S�|G�	@��u�kRLU�������8�㍂�W�#pO!��sk{�lp�ȋwߊJ0A/��'���؈:?�i�*�B�t��|���&黲��C®�s��U��/��7���좩]}<ʶ�rX!d�c2��Ay��FE���P�4i�����$k��y����8{�&��Ď��%���o�*��7XYȪ/E*٭>��M�k�e�\��^@� 7�a4���W&�V��g	�MI2�		�&:��,�o;�&���tGS=o,�^ۑ��¦bk~�9`�!���6��M""xI��ӝ�zQN5�Cj@��&����V3|z�gVl�O
0�:�b¯\t�.	���2��1�k�� ���9��#�"���&Ddr�o�B�?\r�W2���q��
��Y�[^$u�c`JƷ�r ����V"}�9ug���T�Iة��䔹��Ge�(c=W+K��K��$�S���ٺ� P%NEG�ks2HB���n.D�{��{FF��a��l}��E�$�eqbSױ�bz��w->�Q���XlxVHYEB    aa52    13d0���6��]3Ng?����������4��"J�QS�
OynUK<U%>�-����P{����a�{	��C)^����]S?JQ�|���Z�w/�D̃��蜊<˰��N>�ǣ�;)�Uf����;��c�8	�&�M��fkɿ�/��M�
���vXЃ9v�7��@\?��
�ډՇP�4�_��^U�A� �#��%�l4�U>	Z��ޞ�c��&"�D��&	�E/ɥ}9:��w�@�ɥ�KF�[|��^�f֪���:%i�^zi%}��`c܍'�}�i�Den�q): �o�5ё���>��9
����I��I�yD�l�>蟹��Q2��2��ƿ�в%jF�*�-�~|���Y��E��\Nv~w�5��z3w��x8�˳D�]����TD�KwĎ��GZ-�n�0`jY�rxӣ���reJ=�����\��Y̓�.�� X'��g�����5·b����V^`}9L>�� �feo�F�9��Nu�_�-hP�	�0��pk�T�hJ�i�2')���}X}a��_�0/3�O��V���9�!������91��T�FvB�0ń���f�0m<{��]��Q�!+Op].Q�#Ō�/�]��֑��yJ)�h��mr_
l"�\L,�1��Z��X�G(̘����,�buk�]�:��	�%"�ѓg`h�<� ��Zkֳvs4]����ڜ�H�76kq</�͆���"�1�h�X-�º�U|h������DM�����N	��e)腰�W��q�
���`:���1� ��Vm2j�> �����ќ
��E ��_�ξ�t�kԡ�h�#��/������I�^4�Ƿ�ebk?�5H�����t�lU��/"�
���m�QM�a��.�'��&ȅ)Hny���qyU�1uXQ��mo�y�����|�2��=��t�Bm��c�y�wJ���33 S�i��$3�z��ް�Y �wܤ<[���4�4G�R�,�3����bI�� ���Nݞ1c�W�T���'%�q9�A�3���U����/l��E���N8�i��l��p�`�Qez�u�����n��C�D��,��{���M"Ѿ��~M��(a<�-n�I��i)�xx�W����;�pd�|��G�el���"�dq��P���ޑľ
��v�B�����E����I�٨.{����0Q��i���S׋?�*��q��˥�#��0{�V�FL\�k��k�����W���Z}�&�Bl�jy?_k#Lf���q��Km��+��J���G�����E/_A����#��&ߡ�v�4��������('�s)���E�K<�� �����B���8�c}�Ch嘻�o)�Zq��[%}�7Ky�<m�qqV"~a��I�3��"��k����rK�y=%�ۈ͗L���M�@!�]�5]�+�yD������>�c�ƽ�us�ųf�?�)U}��&�v5M�i�w����3>���(���	�g����r��ɜ����@S)�u�߁�yS�^�C6���pXb8"�������SpHD!��b��˻��^��=���n����f��#��X���lZu�耖�'gGz���J����@SNH�4��=�K���t��OJ�*,"�iG ����Ho3�&&���~�w˘|M��3@-�=3"��Ay��d�]��vx��a���cx�^hb�3��_F��TB 6�AQ�HuMt�җ�!jU�P	1+�1w^��=ʬ���V!��_�8� ݪY�k��=1|��{��^Z��5&=h�%AkÑ��o~�
���6�Oho ���;����k�Ւ�8I��O�o\��
I����$f� ��w]���s�3	
���/B�_D�Og���\N:/u��L��SW�{a*���3_J�~lH�F��1N�
�4�*	��G�o��p��� wtGvA5�H�w�C��*�@~q�,J���"���H�8�]���mS��l�䂜��>0y-ȟ���4���E����ˍ�u}�TL:�;�:��#�$#�hd���o��Cl�3s�W�ģa�6�\-Z;��-��E���ր������zj`�������&�E���|o�?�J���.��Ȫ�[�≎j�h��^�ӌ��:,�Te,�3`�e[��0��d�>�&�?��糝�p`�h�Cc�����Q�K)�˗�^16
'�
WƜ�/R�utK�����=o�y�a-MM��h?��.񈢘�*_y��b�u[ ���;�d{\���ϔd� �k��B�H�����,v9fC
�S����߈N�I�xa\�?�.k71}��ܣ86MW�z�p�S�!���[�O�6ʔ�cW�k�c�)&7�)����J�i���E�#�:��Q������=�:�K�'��a*2KZ%�|��x���g��@9S{z��5ZnRO2�ډh���̴�&�!�<���C��ׇ+���+{�h�	���6�'Y���0J�.��2�X�%H�g�"�B���H�(��B�&`��1�����񔩁�mG���� uя �La6�'�M�1��Z�h�e�8%�,��,2q�yPlezD�n\���ɿx���G�v)�,�����xs
K(�W{�W�-�UI�sL���d�w���mc�d.E�����M���z�egR��v!/*(7R�����X7k�L"�L����55��[��`:��Yh�F�G���u�/���:i����^f��-|�+�ɜ��8w[1�T&w�2&n��L��{8��0�Ա�
�������;�#Ac]%p��P��讧#�����dA�u��jV��Wݓ�,�S���o�I;�e�6m^��:��f\t=*e�M������U�_�c�N�����9���6�+��Wxma�p���=^�ʔMy�Po���o;r��[���R��:c�ϴ}	7@Q��V��?DFŗq\���kj�8�l�A�]��0h���߱�6��`A5�2'? -.��	"�� ��{
�&�\����dP�I���&�9�
 |CSM�V��y����4�J����wb%���iu��k<�(�|	#xZ���y,!ڏU�ܱ`U?"�~F������e[uh��O����` ��,�5-��u��v�%Ҷ��JOfcvܓ��ɸ�����V�on|'H�av
r�Z�b��:�#��؃T�xXk�E�H���6L3�Ge>Jײ[�"hh1����K칊�cG�z
IFaf:�l�;'9���aA��G���Ųe��7'9L�i��a��D�86F���V���ņ�����;�x����΄�D����G�<��0Pt��[ǲ? �5�m�H@�)"�J\׽E��)����`Z͋���"O�y	狟n���Iu���'m����(��)�G��@���(�_�����a"�'���b8NT���?��Ƣ��Ւ����ģ���f���[<M�1��t,�`����o�_&���ю�(8V?y�z/���~y?/��U���p�}%+6�ʴF�=��m$��(��Ҡ����\���{��)�&�w[�����i���r���=v�>�B����U}��녈����A����u!��0
ȅ�u�\֟6}�P')7�Z?OP��s�&V���4:���E#]�ְ����C�0a������n��ա��<���eK)�6]��/�L%��"�TJf�ʚ���y������O�mKߤӀp�@A�2����5��r��2�tҋ�G@Q1`�R�k��K6�*���=Yg�q>?p�>}�'J1��(V��O;�`'��"(?��ƞ<̄e�-��f�E��F��]Kne3C���g�ly}3i�nm��XVN�-k�Ih1�I$I���mrP%V��Zʮ_!d:f�o����E8���T�g�Ay�7�Y�76���`x۬殤 ®ܵ�vǤC�m���إT����{ث�~Y���s9@��0"'Ζ��||8"<���fȏ?K��,����w�VÊLYE���AIt���b2��q���uC�=�tf#�#���g���i�,�y-Ӆ9�ō�i� e��!�ND�aC  ��-�Ք��隠D�}�En�#�zؾ�f	�,�W9c}������쵟�^e&����+��Sa?&sz
�����p�(���0� �~��0�[;P���)RRj���	]������g��(~��d��ӌ)�/�����f.���sN�Ъ����h�9��yl��V��\?�hm�\���T��_���B�U�DlӢAiC��B�����7���Q�����2�*-���~,Z�L�I�jv�_�S"<�\�.��^�<J�e�o��i%ۡ��3���]�0J��w����HG{�1j�B�u�uW�O��ݽ����gܢ�����kh�=<qˇP�d�;*����MT������1�w��P]����G�� ��"���n�q�%FV�P��M�\�vp.�U�\�L.͜㸳=�2��Ĵ���߾�F���e�j"�b�$4�Șx�eyӥ(�2�^��Kv>��p%��!��/v{!�5[oj���a.�3w%͝'����şd�5���+Y@1j���Qvv�	�T��.Nz�!b,ZoE�d�����;�SL���T��6�'����)���)0hi��*y7L�݀�8a�.q�~/����_E�b�e;��Eڗ���G��"��'�,*�;lE\�E�����m��Rsև�:݌��Ȣ9��}vsH#9�X��D�x�1w�߉��x�zo��
e_�����	"�=5&�᡿*S�Nf��n��)m��rZ����T��&��5�czԥ- eD��������#�f����h����/��A(�J/)B7G��e���hXQ"?��^�ǝ�3�"M-~f��q��f�Л��d�1��e�QIs�I�z����	�GK�ʓ#��bp� �Ȫ�)Oid�����[��f,�X�[.َ�7��I\��$�㦰�{�R