XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P~J�`p|L�I!L%G�����;��r?��I����y!k��X���L�ls�2'�Ј�|����ѭ-�X�G��<ˉ	�F&�KP�U��E>:E�u���1�yA<����|E<ڨ�z4�ئ\����w0��rJ;^?@��8�!0~h��2*`�7H{��;m����p�)z�wKl&0�(T���q1���zs�e��Y��(��?.�����$XZ�����6�*_0�N$Od~V]��(-������<�at&��#B�)N֛?�_	��T8�}N�c��s=#[q���Oe�V'��*M_z%�Zu}��ь'���z2�]�2__��ޮ����00;5����5UC���ʑ�]< �<�b�� ����R�J��7Г��!6R`�m�t3���b�R$��.�9��G��,�D]�����Y��3�봂��1�w��Wr>�
zd�jW�'o��i�䅤��I�f+w�uBۿcob��X���OV���f�{�$
���'�k>U�dY7��F�J>G¡�L�$e�㢅���P�n�~�Y��;�yq~���۳m,�s���2�q)�p��tf&�_�
�A��$���"�NZV�(B���r�/���eޜwM�4�����2)��s���>�t	y�X��F���ǿ����L�/aq�k޸��6'�F�-�@})$��U�I���QP�vjuS�;3���pF� ^x��U�&�B�d�ݜ�v�t��ˣA��Z���-����y��XlxVHYEB    fa00    28c0,0O����!�����)HY��x��)v]�|�/C:�ߠ�)��jzo��'u$O������Q��Zؓ{�3C�+�g���Y���P����9ƻ<�r��p�Lj�W�@�l�f-��'�9�v���[Ɲ��$ķ�����V�N���i��r��f���R9�t:����p9�hl�@(,#��eP�M�٢��,(�ww褏�Kz�W�>��P�B�l��57�ʉ��d��]��qź�rY�e�T~%�oEF, �q�`���,b�#-���/����f(*�<8r�uȤ#,!*�������5�a�?������c��{��&m@:nj��Q,BW��,s�M�dgg��h��C�uc��q�
� �a*#t5�e���=���Ʊp!�m_nGf�0Ad��^;��o�A'�*A_)(D��γ���p���c�^�v���QDŏ�,I�����MgV������X�/��p�x�?YY%����X��<C�D���B�Yó��T)ΐXd1h�,VTS����4��jQS�w �h4	S���q�f9����, �����uӔ���D��
L��ӎw�:�����ᑯm&����ݹd1g��/� �������I��h���$E��M��2v�2�Bʹ�`�L���qq�qYI+�,�.��WN��-$�������n������gЅ.0hٗz�2p̯ �2�d����z�&NSBn�O#/L�\:�Zw�A0��y.)BW�!�N���۱�L H�C��@�62}�}�����7���RV�0\w�+�ߟ�2_"%����r����2m�
J�\=�Q��Y�g�͜���N�nMz*�c��(8��7b�e)��@j����ӷ��i�D��R@#`�#�MXˬ|1��O��Tt�����v%u���4�(����^�=��g�~m�7���(����o;ݻ��T��"m�G���i���@������Y��԰^��+?�_ՠ���Yb��d3�!�[�BA�=Vd���N�aP�sdȜ�I�t�S�e�2(����pB���*�%�;z�
���~���2���{�G��"�q>�Cr:������<�V.`=j�KǺ�J��)�N�c$	F-���]�{S�B��2�ʹ������J;�ql'�
y|j�}����I����?�$r���7���j��RUP��P����r:��JB��0���L6��$/�� !߃3v��B�Ë�����o�w�����#�ß�W��o�Sx������m�z��K��q`��K�hq�}%ĕ2��a�v�@Gs�������I_跇��`�P��W��Z�H�`�&b9ǈ��L�6�m8*C"J�6��D�Qۍ�oB��Q!�N[�N��U�����ɳg��U/�{���"Y���<O�Md>����:�/�,L
�+u�x�yK�v�j/��kG�?�� �=̔�YU�VW~�9��!�阢��]�y�����R�[��r�M��9x^�X�3��>�Fa�hÈ��0��o_�IQ<�����;-��:�y
AVb�75�ύ%3J�>L)	�0�Z@s�0���,���b���Af�!��CW�>�}�/ +�<c^�Ԩ���P[o�\�	�%�HC�'�C�t;d6-�n����Om � ���֦�V�D"wa:�^ߣ�|5���������.���m-*+��p���`���s����B��<���X�Z5;Žp���mp�S���t�g:z�|#F(���U���<�H�LmX6���y��e���bP��`�վW��`M�I��ė~~V��k��=�pϢ0��KZ�!��r�ʍu�#*e_��w< Y���5�(�������ӗ����ug�, ��r��q��B���IR���Ć�
��uv\�_�s(o.�l1�O7��v52��/�<��DnK*hE����!Eyj�A��U�e.f��WG5U�A��l�*�`yȝjsc>"x��BU��ސ �W &�"(�7���}����9s�w	~SV�g����޹!m)���᯽�6�U��'7�5�/�2��
Q��I3o�o]Y�����3���3��r��p��I��U|�����	�T��Wr&�X1To��ʆ���ɟ -� ��9���bF�[�|��i)�Y�a���U�]�OW]o�	��X��h�9s<6�X��OE��|�^�B':�w�L�2%#����r�����-c����V�CfQד���E6�SM��*2�}��������ؓ��[� ����'��@�����C�~ǡ��]ͻ�	���Vl�r|�
3��qXt����h4�?z،g���m,;�ZP��u��sy�-�"TEu��N�m�'5�BrBi�í�
�յЬ@L���dp��apG��qՙ��պ�e�"��G���x
u5ZUd'���Г,�����{�+��I���7���f�8d��y� �Y�#1�;�s[UU�s�΁=�FO/c��V4D����ܯ�"�V�Xw�Q�����wX����V ���|bR�D�c�!���L����B4E���Ht��x�C,�'�ZW�\���A��Kf' ����J�g���1����ʠp��$� &m��X2���vKܯ5s�=d�	�4�����t�f�R��N�]UQ����g��\^�����v�P���Q���`e�u-A�<A���!!5wAf_u����S.��2Ԕ� ?n�M�J=�'�r��jo������֏`�o��l�ɒ�06sI�1YխAa&���o�%�̞�7�)|k�/��H���P�&ad`3��625�չ8���S�����1�{ϒz�"����.���HW�l����]�����ӄF ��4[�ڀ�y��+��XR�D����ދ�"/��������vF�t��1gs쁢�@��7�\D�p�o��]��]I�e�=���x�1e��9vh�np@YJO��'�{���)5�.i���fH?���aqp�|Gx��|5��]���;���){z���ћ�
.��{�ݢ�V�~5ܢ`2C/��I+����d�r���Ώ�'��ܸt]��t��2�n�bx B��Yq�M���a��}p.m8�^*q�a��PO�%�Yer�ng�0!�]Cf߬D��ܕ60z���y��_I�%��B��J1R��^Mt���4K~�g�Vl����ol��<���w<�k��o�es�����%��j`�g y��U��s))�j�J����'�S*����bC��aQJ���נ	���o��ધ�o��:@a_�(���N�O��W�tJ��|o��1���~�w+���+����W5��T�ȝ��ކQ�;�O�Ɩ ��6�l�u�a��	z�����-���W;�����i3]��	�í|Ng1]�tU�a��-�c�y���I��g/d�"\���U�5t��lZ%e&���T4_Zx�ݸ�<E�3�ϯ`-[^d�n�~'��8�ޱE��e?����!�哀`88�Y���U��AV7贪�Y)�[ 3coK��[%w%j����"9�$B'yW4$��,p��LQR���7){ߜ�Y)��?[�
�E�H����F@�kO��}R"xr�=�4����_$����i:GO�m���|����Zd;om��%Oɦ�|1a��K�Y��;���Q��G��Y���ϕ�?����N�k�,��jv���'3O���n��U�>/���P�F ��z�b?�8Zݧ����dD��S�~�4f2��`�@��%�����������NG?�U{\(�X�K��f��OL���b����:9�OPAQ9�dHLo����x?_l�I����$$�A�\'iVE���V���kbv&Qq�����V��Q�sƜT>�>j��M(�'[���%�Y��!�TY֧�\�m,o���3�.g5۴�����p�@��M�:�%&
쥝�;� F#'��;��68�`Y=�n�7AQ�^�_d��L�����\Q���Ôa�=��划]���G@s��*'�0����'���%,�F�iT-�1�,r I<e�U��(�Ϡ;�����N;��2�ɦ ���XsQ�j?�].�xK��Oר(ij`����27:ډ�B�D��WF�]�����U4��h�*�`(k�d�m=܅�̇ ˺>�nJ����:�޺%�z5�F���B��0ƅ��7�f�� w��P�V\}Çsu �� {�'Yt�!��o���M���O#"�x��_]H¿�鏹��������^!����4,3&�uK7p�ha�{ǭ���à����<p�<Nνv�%�,�H�+:^�<�`�\ot���#м��~��b"Cs�ry�#�V�S�E�5����N������K3��8��4��a9(��L���X��)AF��.�bj�=�F��4M󴔩���r`)�ďW�zcÛ�R:WE`BFzG����������(?��(S��w(�P_��?�ާ�f��x����:����`��^L/����QB}V�*K+��L�O[ �oב��"�8)�Or_ٍ2ݯQ,��?��bC���Fy4�g��Xj��<Z'�B��=� c�	L�t8��!��dA右�Vu!\�[�w��0,�r3Z�'}�\/�P�dB����^��ҦB1�Gv*R�w��]
<èJ56��G�WS�_��wJ��BF��'��d����oAB�i�;wM����/	�A�1Tx��.�z�D??��+[
V0��X�)�ﻉ�<�; �	��I��U��ב�����8w�60���e\�P_��(ѯ���(em$k|Y�'���+5L���<�(�oS��Ŏ�R8�=��+���N���-�h���� . ���b���h�"���8�QT�O�m6œJ�9�y�)bB6~��d����:�S����7�xO-�K���N�b?�B9G�,��2��� �؂>�5~y	��xa�9�'ya�e��:,���T�0vI��n$0�TOp�ߟ�W"��t�7N��:�Q;�eU������]���A�Дt�.�����#�I�Z;�9�O���)S���W'��t�0]N·���Rכ��juI����w�·p�5V�P��#TE�����7a�'��!~^��+D��6W��{Y��c�����H�R5J9 ��hX쏁/�ѥ�Fk5	���s6������]�Z��O{�Sz�7��(�맪�P����bG�4���̕e7�l{a�M��e0�TX����^��wJ��z=`�/`��D�)T�7���
%���Rd�Yi�f�I�;_P�$�Tv�T�6�zw$�0�(�J���X�"����SK���i܇���c}��4ө�2�����F�{��YG�N��/H�ٰ%\�P6Ȏ��RYN���z�<�+����z�����Ӆ��%��ܴL)����B7��!��v�f�)O�&e)��g\[6Ϡ��Z�8oT�0��X� �>�;����`@���3���c�8e1�(����$��o���p���jY�\N��Z��q[�C�B�N��FQ��S%�;	C&�^@��*n�f��I��g��+MΪSx}�����6P�rS��3�x���m��6G#�y����BY� 9y>U��<���Sƌ"A]o*(xX-z5D��Y��&_��G�T/��ya��d�1�Y�c	�hG�Ny:��� �kLp��ƽ`5���K��ך�I�L�0f�J?�"����h�m3��l��xs���^!Y�NΉ��r �.�=�})$U���<cY*HgU�l[��3@���U��S���~^�T2��_��$�`H@@35�L2J�N�0�@Mc�i���j]���%.B�&G�����#�}��f��;�vo���N�6<�>{/�e�QP�yw�8NBc� �|d�<Z��M��t�'y�k[\ik6NclEuI��vz��ݳ:��d�~e	;L���;O�9`�L�ϫ\�*v��e���ߣW{o(���z;e0C��&r���?��S)�4�q\J(\`k�1W��0��m4�oβ���v�t��;�a}�v(�������t�u�AS#P��Rc��
��,�f�Vy��W!�h�CJ�d5X]�X�����M#C7�SY��N8�Tͤqd?5}��7���,������Fm��!�s�"+���3F��U�"�/��5C!���2<Cu��k�YB��� ��(.\�/���T#xM �y�S���n�L|��e=�.�]#��,4s�?wE�����aVC���9nj�-͠^��Qi�z����a�1��1����a�I�tm� a��*W&�����Q�$ϓ�R(�^� U5���{�r�|7�Q�Cj��Ŗ��*_I�������b������؝1U�����t��&�hB�N��j�<μU)�&���Q����nXMKqvEo��4�K��P�͏un�.��$ە/b%/�
eB�m�1"j1'F]��N�=����!��C�ݯ��>0�
b�XP��ez^�^�kn�|� mVT���GH#�0,RR�VFaQ�眨��1�K�W�_���y��]�L���x!��P���`����b9)��&�fn��Z������Ft����yD���2�_�6U��{b�}������#I���)�m���2\`����4��+��k�A	��d�7E�y�: �`��U��>)��s4�.<Ŀ�	�^U'���Z��*����>��_�קW��I�������LN�x����=ŷ���K�)D���zWm�{)3�zW��O�hn����z�`=��ͱO4h�_�C0��`�-F0�	��R�./����9M���|�}p&�]�蕂���sBC[���2�Q�)��0�	��$�Op2�sE�2�mDF�ə v�:���]��q)�6����E��x���b5�{+ʧ��<�R5�֬�g�!Λ�"�&SRe�=����=��%P�>�J�4�U��h2���Cǣ$���čqK�!�ި�l�� �� �3Qiʣ�/?�4�!����<� P�O��:�
q����6L��7��h�b�e���}�.��1���5�Z.8$����ܠ	-%�/Cn�cDu�߰BE2����%�i�4����)�$%(")�@�߅�l0��>�\]]���v�لW���� V/6���T���{��F�@0^D�DO2�_ژ�;Q��U%}$X�u��f�����Dm������,��n6'�-|-�s�
���VX��EP�,��ڡ��+Ƹ�v
i�Z�D����S�QKLȅ���∮�p���76 ���m��A���>��1Mf�X:}�Z!���f��+~!�0����J�f�1~�
5�;�_�����x7�'���� l����:�v�
�G�R�J�je� }ɽ���߫r�-5�v��!o?T:2��VE�I��{8\��y*��.���cl		��>9�@���hm�C�خ���fk��.8��4^���L���H��a��[�1>�O������������?RFPum������ ��>�qޠ����jH]���e�J ��(XjT(��U 7�2ʫo@����`��0���g����Y�[��@��0@��a�+���`Z��J64wx1&�G�0!�dk�[e2����9	h�屮A�K�=��8	�Q�?�+����n��g}�R����F���M����幃`7�x}�m�s��HI�T�8B��S�����?�Ma���ϘB3�ޝ�hR������J*��kPiq,۬������h�7V��!/��̢�:c>Ƀ8�L7̭�B~N�MnwO�)p������A�j��P(mO鮬=��l�.�2.��A�,}#�T8�DX�Wf����{��՚���:r�鞈��AմV��$`W3�ӱ�xڛE`�y�h�ެ�lH?��!(ul�iJ8�W|�/Ŵ�i��W�טN|�}}��B������x~Be������P5$��$.��:L	x/0�d�՗L��V���s�%��B{\ �"PU��2�͕g@t!�A�t��ŵ97N��;�W�:�"	UEx	q�m�c�`W�P/����9o^~�p�M:��P�*+��4j�_�&���� 3�s�����r�q:������/zU���KB�Y��e�5['�'�}DI��J�[P���N	���l������	.��
����O��1zn�����^b�4X�Ȗ7���w�Yc��\�"'_����+�6L���n8^O�^��`��:I�SeB?�u�P�k᷎F��ס�j�"�{��l�f���,�wXH{}���h�Y���c	+�x���q�}n��0"�K�Y"�l8�@r+G��'���:(�xx?Dc=/ �baR��2����w�~��	b�����E�NQ��d�VU� t��k$/���=�Ѱ�����Ԇb���<0o��r�k������b��C^#a�ʡ4u�U��%��}��<�Cs����o��NQ�@hB̒Ib���C�*~�Q®M.o�,�M-5]ʋS��} GdM���3��臹��)ų�l�Mh	�� �`?f���0��'KX�����Je2U�А-��tMs>t~��@�;y]M:�<&�'>�t���ݡ�a���|%�-��@9�����o`�H?��&��B�%�E:`&Jpd�}�ENa_���(�d��{o��*��A�&tB���55�;ſg��*8�F
�A_�d�q669%G�n�q�s�j��Co� �E%b�m�"�H�����o��#���ֳ�D�T��QQ��k�@�y��r��>THm�- D�:�-q���:g	iu.~N8(Nq�4�
Ŀ���K	�x�!e�4~��f�,a���Tb�{:�J�$��n��inJ��2������g7�v�m��E��d2b��C����v���~�������'o+���r�_����.@����6Ęo��J'�I�b!I�ne���4[��#�h`��b2������Mj�W���u�� ����Oq9&.~G^��%��A��Qo�����EMb�KZ��縪4���f�K��J��9�a@Z����)W���/�x7r(��?jˆ`���[|�	Ĩȥ���1�����@1��d��;uF���}�e��@܋~\{��i�����~�,����(YL�����j�m���ɥ�M�+y�_��ZuD����\��(?�Ǻ��:4thf+\���G��?\�N����G�2���n��JM̞R�S���)�j?��Y���6��?����k>��*�N�w��Z�3�8����4��j��""��Gp�31�bh�/V3�Q�B�~��V���'e�/x�a"�\s�'
^
��Qh�zE	 d�HENC�>�֗ �R&W��02���>�7`��E/�������f>K�N(�`*�e^��4Q�ƻ�'k�;���	@pP[��<�}�#����wX��,�Q��I���>j-�Ɇ>,�C�)=g{��v�|\BF��r�����.ٝ��{��X>�ɦ?�ݩ����w�a�`sm�0
� �L�+�aܜ	a�X��I��>�����+�0�����I��6@@R���PM~�����G�B�#p�h����c�/��4y��^Z��8�,|���[B!���=����F��̲,�;��'����?�� >����f��oך@IB�7�e-���}4��}����v�ܘW����[5�P�(V�@駏�{��~Sj�o�gǍ*t�nL��Ǐ�N^�<	B���8ٔ�G�p�S�[���I�o�J֮-1e�t�p:���s�?�Bb���;|A+=��	���|��{c���v�}鐕�ڱC�QtXpoB_�ϒӏ���'��'�{I���G?�>=��/W��n�Љ�x�2 �ڍ|��~cK,Ŗ/�b�n���Zp+�S�\��"fN	L���A�e�!��@o�/q�5W+��a� �]�@p���T���`�S�a.�g/f�Dj��8��p���&d
��GU�;*���M����L��_��B��K�������eX�	�o�nU�l��1E�ά����W��q�J=�#]���~|؏9�q�h�y�f��z��S%;�& ��jՂ~��<C��ӌ�r4RwW��0��i��=�	%]t3�u�m�xDY���A/L&���X���Y����,�H�H�ܥ��Pļ�ń���1��*yс�����<��%yC��!�[K1C������nl��V���o����!��h�XlxVHYEB     896     280$Ш%G$�K��Ü0@�9pZ"^�y��LyQ��r˨(�Z��vlo+�\�/.�=�C���'�4��wT��
׬�cf��ij p���+��G	�<<�^4jt]�{o0���
?��>�ib�MOB���B�`�5���Ġ3�P8[��s��]���>;Y`�Ŀ{M�ۤ<Ԁ��İ��@�7/���:�	wx��7�u�Ds����z = .č�\���1D�]�6t���-�>���]�9�q6*�9��K���e�����F��>5����ؓ{��#;~�7�X��k%v��}�u��<����T�45��L�9̵/M��N.�HS�k�ME�5ژ�s�k��勩:~N����ڱm]�k!�ĠnH/C�B�S	� Ϳx�'$�N(7�������a%6ڳ���iY�!6�������GnF"���%;�n�A���k**PL���T�����1���d���J�����<����\1kS��#�Ϛĺ�S��k�Ѷ�=[��wƴO���"���߃Ͼ+�v�[�>�+�3n0��K��rp��(X�G%��!��4���V�V��'�.�gh��i�O����K��LU��(�\�d�q6�&� Й��\[��]/3]z �