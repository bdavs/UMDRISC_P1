XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9�v�2�9k� �݆	��S��\:M_җ�I`ma �� ��"�*�O��f�ei���t���՞Z��`����bP�B����<���s��D.�Xs��Gag������vj��]�|��� ��n�XՊ^���Z��@@>� 5�xAZ�_��N�ȳ��'PH�� F�A����r<(�o_|[����	hJ�L������M��0+N`�s��+���?��gGy?V�o���6�SIkYU�����t���<c,���w�T޹��%�UHo�a���t���S���L؋�-�C������M�Kn�)�4x��w� k�C����H-?p�"��,�Ruw�Z���W�Ea�=����7o$9d�T�,xG?
�� �i�x-\�������� tp_7��C�"�[RD~�>�l�uW!CW�T���=F�
�T�B�K3��h`n[u�39�����/&6���W	�z�`+7�AԷ�����=���4Jx!���~�iOӍ &r��cw�z�. >�����E�����<#�2}ٙ,T���7!�>e�Q��F�a�E��FԼh\�3������2����q�$�2r;��~1�T+�9t$���O��Ic�z� �Q�b yצZRĨϘ�edF�Q�xxK��b��Or��[V'�qζ�Pw�r���q2uO��l ���Cԩ}�0�T�v�+t� ���y~�6�]��Z�~r��r��!�is�<�hM5XlxVHYEB    56d2    12a0�6|y�\a�%��OnU�.,��D�i��V�	�W�c�3�B�x��TmX�6o
��I����G�O����䮵@������4��"e���A�=`?�����%R����D��^;p]@Xz�K�]��|�ǲT�<#���O�-�lU,Q�;�8b�p�P"'��^�b L]E��_�]�̤^��O�� !r�M�j{%�
�QL�Úω����D��B�J�>����-�Մ����	�X��"�⩣)6
�φ�7�A�����4
�K�XmsA��M@�������ƭ��}	o��xor�9ʚV��x���J��u�'�kN+��./U��V����  ��_����lWY8B�~�dXh�cˣU�w���P�"���>�Q�s;Q�/�0s�u�x9[�cګEp>k���>;a�I�иE)�FP�&�������W١)��p����m`�Ń#�������G�bFj��,��C,D9{������)Q�
�Y/nq���%���+�L{��]�8R2
u�|��M��Qz����g��Z�ު�Y�/ �M�D���bD-�|�E,����4BPu(��1��]t8_��2�P��Tk�V,�89Z�:��N���rR�'
��@��r�ct#�(���c�����/�;<6Wg25����U�v�"�͒��\���/E��w �%o���m��vE:||�h&/Ě�F+�xx����O.��u�o�MC��'{h��r�n��0L�q���%h�)���t�R�C ����*�0����6��b��f*=Zu��|2?e�j��P]��� ��[[��K�ŵ�;L4>d�a'{Ef޲�a�c���I�����Ǚgݱmo±���䤸��b���^X���)}�'��gA�A����ȍ4q��*�N�Ǯ��Y�@�mV�I�U��J*ս@����"�0D[q]����<@ڈ�$�>,?��+C�O���3l���{x�>ɢY�H}#�d�)�^� e�����N��-�)5��JV:CPl=�.�K�=	h; �%F�E����Ny1R�^k��~���{}bP��'�]��\#R�|R�ZK����-�7��눣c4��.�[�a�ټh��w6d�P�w
��ΤѺ�m��B���-�p�֮�U�!Ř:4a^: �̰�}��V-���a�0���49\/�__o�е{N&�FV+U�2���^_N�͡4��@v�&�@��@��sC/2i
��C��7��h����~������g���\lLrj�/^��7]��d�6��7d��k��#���C�[��Z�ܫ�,��|�]�wgY�\��`�#Vo덿��)�I*��o�ؿ[W$���KNh�G�3�:��fϘ-r����z����{�������F�������7��%B�F+������!,���JtR�|�B�aJ�3��z�D	��9`�"C�<V���+��.	��.kr�1H&|Tl��&"m�j�T�XR9b[ņ,� �Zo���:L>)���滂$ND��vF�)9xU�
��%�]�a���RL��r+�g��%ت����^��}������}����09;$Ξ��?T��ܚ�Pꜷ�/t~bX6ڙ/�o�/e�+���ї�Bk$�Γh��8��a�u!�I�Vj�QF7AA@����(u���q2]�������mUBp��e����y��a[�3�m�ܡϻ}	����������	ذ@3h��1����Ͻ���(&h@�"���4>���f�� �&���Z�ArJ�u��[�"Zi�,��N�ǿ�/j#�Yjg��+��t��.�2޴�YY�wռ��|7Si&�� �=��.m��;G�m�ҿgUT�x���W���[�Bi}?ĥf1o�����-����A�H��Z8���7f�2���&���^*f��Y�d�K�*�k�k_�$D Z0�+N��2¯V��3�4�5�g,�5�:�2M�t����r�M|TM ҵ��Y�<#��Dǔ���'���C0s?q�L�9��Imǆke�K�o�U�4.����5.��S���R��'�����{�>��y�uyƌX�O�A\�ޖ��"a�l��Pck(�*c}
��j��k�A����֧/�8�NkJ�$S�����U���r��|e�N�Bb�=�9?u'Eָr Prt��Z�$5���䨛��v������F"�=�'ߌ0&n�j�H���l2o���ߺ��)v��>	��*��h��y�l{�5�e���Zy�O���&��
6�����3l�k���I�[��3�%��˨���4�p�u	��7�]�Ś!��)��mV�=+�n�<�y��G���O��T\��E^/vu�5ߞ��3���أЖ��r���J��Sی��y�k}�qx�-���<�.����Q�3<|�IH�60��^2�O�,�N�����~�;����#I��>��/w�x�>����	:�f�� n3:���S�H�Ӂ��`�qd�:|��Ѥ�:2J0�V� ��9�����LA�����Z=��Y»�,����/��+�u�2�@ϋ�AG�&�,��I��~+�����U���?�S�:�=�T�)҅*��TXZ+OPsͻ_]�)S�\�M'C�c�*�CB�b�o��ⷥ��f[���T����e<�Ai��U)��������wۯ���|Q����W�P�'�dm�9$Y�T�g��%=��[~Y�ț�H�2ʞ߯a�ʋ��a3"��t>�0���C(a�֫4`��iZ��2�p׫�i!��	3�f&��A�Bv�x��zua�,0_�Y�� �)��h~��Ҏ]���5���ɢD�o���Dq'(��������k���!�Ӫ=訡�J��@;쎤+֙��K��8�	�Rf��^�j�},�Ϗ<�:�cţ��w��Xq;���W�:cj ~�C@�(��eÂ�2d��*�=nꄼ�c�ΆU����Ǜ o6���z�1T$V�#�8!H��Y�|s8���o�)I���du��߄�I�3�	B)(�n����M^$��v[���I��Az���k(��Ќ����i�7��84U�.5�7�p�T�"d�.�E�E#���FR���DHc��9j	�x��~_h���,�ͤ���y�74i�%,/ۈQT~�zpqR���q���g����)��	��KL�����}��a� ��沾���ϧ�ܘx�yօ������M�F�j��Ϭ�!��� [�j�ϒW '���֓H�7_�� &�T�/��KD3FM�&�Y?FY�L��j�4��z����!���,�L�,�Nv7�s����}z��ې���S�Vu�"R1�jޙ�$���ʜ7�V�$�3�7{����$�W,J���6[�U���(�����@����[�g�p��jĥ����]��N�_q ��#���YO�ݠ-����пZ���"b���
'��`���4�nd�")��+���I})��\���R��Hr�qI��<Р:��`8��)����ƨ3o/��͘�� ᰅY���y`I�����u��¿�, �����g<.����):�l��M_̳�|�c�v�X��gɒ���1	��Oc�;��Y_�/����A֮!@�v�C(�B�:�#\�Y��͸�������֊A�~���J����G��L��Xͻ��$r�(��s�c���i؋�c�&�
kDy>��Ci7��$~�}���+�r�������(�Ʃ9'��A�O4o��C�i0��nL�#�0��+�:^$�ry�Rts5���K�C��C�+��Xw���c��� �F;�!ZGz=����H/a���H���ŭf�0��>�_����vxd32!�֥��.��!��Ѿ��jox DLNV~�O���!Z�=�I��=ci���Ld�6kn#;8tS����HI��;�n�|��&�%���2`�ْ�`�j2,��NC�+A\���8*���B��t4� #��.�!~ǲ2�&��$ߩ����-V��I�~ŋ�\ď���LPAL12����%r�ž��wp�7��|�m�^%���S�w>�ԧ��X��%CJ P�\(@��=����`~$��Q
���>�l�%��ڰ���m�I�����d��̦�QE0U���ĮGP�!Z��Ex�)�)�t�&O�s�PW�ʊ�Ч�7˲p�TɌ!9���~[�wGq���~�J��#^�.�n���y2��(���x(t���\5�1��V%����	f�	��@6C&��$s�j$�~%z����X�@N]��T8��|��]�J��y�r���<uʉV��t轛#���I�%d�����aH��6tv׌�\�+Ar��ƼU�W�O�8��3��o�W����=.Nzl���C©���)"l�����˶��Y��\���9���ww�}���Ҝ�b���J�G�O�$3>�p�=o��:2��/���'|UkD?څ8ɸ	�F���(�m�>�GՕ����r*P�G n0�f�?�k��T㫥G
�_��'G/�ck��c�^�?U�H�񥇨��w����e�����c�	9���xf��}�c�;p;Cƾ�-I=T='�!���1Ϫ^��IB<]���~�r���]��C