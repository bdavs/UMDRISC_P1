XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!�Q.�T%H��b �L�E�)��Ka�U�� ��雀��n�����d�R��6����~��*��?y�ڲlt�b����_F�$�����{p#��Ȁ>ʺR�0z�dO�����W���8|x
����k�R5@����}Ǆ!.I�4��Am:��|T��Ʒ�H�B����ϙ#����Z��PS��K�|�ִ�(����eG���b�/� tZ�t�݊�t+%8�oT�������(�"$ͤ������6Ͱ������#���
v�*��b�ӈ%����[�c�����J��e��-���J�p��=�\�%��u@ ʄ�p�k�/�%�Ѹ2d9~ži�s�vuV�7��I3�Q���|�MQ>C��q�h�Sdj��ҀA@��'��>3��{����_0�������o�@�Œ[�7k��W�3p�fq��56��\x6���{pl.%��^^�&`Y�\8�cfY��yˠ���4�,�J�a΅D�<�=�JJU�����!�m�`���E����Yr�py*=���"�^�?;{Fû4W��Z^�nTTD�r��9"!j�p9M2.j!��tj�ݓJ�rE��^���$�*)Z]D	���T�"A�B��[ZB�Jl6�v?W9��3���D<Nﰖ�99�H��%���aQ���s_�'��/4S�-�<���'�	̀����h0���E���3�^N���8a�������t��|Qc2ä�A�/Î��]`\HZZ�˽��a]�'�꘼XlxVHYEB    7744    1780�����8���wt@���S���䟧�
]h<]D��3?'�%1�x��N�}�%],�Afd5fZk��Q�O��1w��~�gj��ȏ6i��zu͈��B�A��5�lT��
�t�U z,0#B�OkXjc�w�e�_�hq��x�S5�g}d�;��#p�! �S����'a����TJ�/��޷�>B�x��j�:���Ƚ�ސ�7V��2���an~+ؗ!/�nfR��	��W�-��ƉJ6��v�z �
��I�u���DU²�'S��<�ҙ�U1��|�{�euR�χ��i��֞�J�\\�ւ�TXnhy���)f>�MH�6I�d� 6�J�	yI�Ȟ�x��ֻ�:*+ե
+��y�m"������F��6�;8�S	K\�|B����@�x�5�l��L} ~d��Ca��r�EA�ɋ'g�5%W���)���}W�����a� �mǟ����?@���p���B���[[�s���T�(��n�ں�`�p)6md�<�ڇ�\P%��Е�#�ȧ�Ld����1���o[r�?����CW"-�ȿ&�7�M:m"ev�F3GuT�Xm��d!�nx��U(:e,>#��D��-�Ʀ��c3���T=��i��mѫƙ&��Դy~��DzYF1T�(�1��:[;�Ly�F�����J�]�eU}�%ZS���Kd�"��G^�돮�2br}�}$��/�%���O[��� d%��*j��:�A1u_�lyE�ά��Ah����[*�!H�+v2��T�����.@%�w�ޚj��YqU���!�fX�g�@q�<��ͣ%��$�%�Hl�D���谨߄H%QK���&4�w�mpzv/��3N���FsX�7�7��@X=���*���:N�#h�,1fe��S���ڤw�p:f@5c�]V[0D���̆�)�6}�V�`���j���ħs�����9��hH���g�Z �0~�C+/���d�S^�^�Z�� ���ˍ��8_�_��Rw�p�
7�2T���\m�S��ƒ	�e��Y��̸ۧ\�׿ݵj'6!;k$��ů������A���`��\�����m�l�ņni  H9p<H�p���G��9j=��{<eo�7m�Q��5����sY���&}H33�yL��x'�J�!,�G[�����(�O[3B��79�)�1�@�^�[*��<) ��9�Xqw���n:U�,�6� O������2z��u����3dX�y�u�	����@�	�i��x>�"��s��6y�#��?�!O��'bk6u쑈aJ��AO�M���K.sp�,�b;3E��g���O`�D�L�S�E�`�V�	&�'�Xx�i�������K��!��'=��~���)(~��}TP��ܐ���&�8z�I�ϗ� ���.��-Z����(b<F�fw:!�H�T��O��i��3�t�vtL�����h�Y0���~alX���-ǉ�ʗ�YHpZ�m7 >f&�P,r��ѕx�Ͽ����+�X��%p�S;�� ��ڞ�i)�@2Ζ;���髐H�r�U��O����5M\�2��h���5�p�g�{Inz��u��w��'ݻZD�-lb�!a�Y-߃^�!/{,�2�!2�Vо���O>��!7���4L5g�Z3���Y�L
Z����]��[PϵD�~�9��������^����p~&.�jCD�<O��)S&�P�}8�
�;@=$�5��(68�M>��=�A7M�E:�q���0󹙸�,�|:�ڹ��'=�ۿ���j�Z�h����/��Z^��◟�c�����9�Xp�w^&.�`Ea~�0HJ�Fg*FY|�FR1����8��=m��>ܶeC��}��W-��!�y���:ͱ�Z�. ���M�p�T�D����w����G��AO%�z1��_1g@ҋC\h�9�v�%��i�%F�m7
Bkؐ��� uD톯Z�Č��>���n})B��E�`ՋU�[�y�b ��F�'����#�{vBi��屼���_K�\��"i�	�H?�i�,�ܤ���Ϲ�k���J/�UMa�۔̥��״}_&�D�3��'~�m*��y��W��-�~<-��e� ��W�H��L�S����8Z��L�	���V�j ��7#1r3�ֺ�b��ę�w�.�/�T�
�gSS�i��ؤ���Ӏ�>F}�RX���<�o�U.2W�R�@���m�u�#K¥2JX�)"�.d\|�+��$�#_��v*u5���V1f����v��J�(p��e.�kM��^M��Ϛ������p���kTa\N�$=�  L���(�{7����	Z$Y̢�<I�����P�+RGW��KiG@k[@n��*Ya{퐭���ٍ4���|@�V�����	C �Od����f����z�Wq<�+��/���7���UQա���R_��ZYg����y�V�·�+�j�;Ch�b�U��J:�/�5c�*��e'�T0z�_Z_w � J��5�J����e�*i�7O>V�l[�J��ҁz�f7�#ٹ���4�yPi�Cg��.�Ņ�4��vN���;4m�x,M�t����&��=�&>8~m����i��t�C�פbIU�0�����\q�H?���ao}v����_XH̄(�6���yN��쉚xE���6wLӰ��s8�Q����	K�z\0p�h@f��e@ʫU���s��@מ'�l��o4L�x=t]�dzs�y�i+�hM�:Ds]���!hՍ�yӌ:u����5�C��J�IB���O~�5�۸.��on*�2c<����7{���6��01�#Dy���� �X�F�~=�_>X���Qjİ�A%��(}��V��y[��������A*ϊ��~�d��9��0C�R�3� �K�%g3��}�J��Q�.d���O�Z�я��s�KZ���Zl�������y��r�948�1ɰP���h� ���b����>P_��"V ��X��XS�W)K���JS�L����Y��Fn�~�\�?;���V$�0�F��o����m�^�U�aճ��@B��;<k�zV�8��q`����6┶w�?��g�o�4�o�?�`�q9�=�S�gp�4󽺌˯�ە?�,SAÖ��`��wZ &y��$8��UoWú�KO	g��L��*w0�*
��6�lL��r}��#UV��gp�*\?O;)�4Dm��?����Qi��%(T���jS`:]��	��6I���o|,�YioOH�G�Î_=S~���$��B�;{G�Q3=}�IZ�Ʋ����=R+)�C����`z�H��jwT�j%��O�W�_k��k�]��*>�m��R��ǝ�` ���U�.���Q[�a�8�-������� �Y�~���A�{ H=pK��o���]���Y�-��[��P³�9�*�4*�`'ڱ-�22)V+�)�ֲ繡���1\���5Z	��QZ:,�}�|K���Rh;�#��U��+��M��G�j�O�o�wx��յSK�4�(��: d�e���4ytK�RJv�,u��^"W���1Ʋ�"�lA��4��8�r_֌�@*J����;j�N%�C��1~/*���?���.|G�V�i,�!��C���.h�a]���\�u�53�p��E��xo��o��:�:������U�y��ǚ��a;��˵�ȴ�U2���G�u؜!/jM@��,��e��z��U��T��F��x���k?�2fž3���X����Q`͕#qz��=׹�"ׇBPZ���	.u�_����Y����H�hvl #�[<.���i4p���l>���9'�1X�E}��d����m���qҢ�f�H ����t�k�P��CՉ���z$-r�����Q�[����|�b䇪���;�:���st'�+��~��C�䕓�� ]�Ў��tP,��j1�d���7q�6�3Ŭ�_�X�C���o.��z�闸���m�8��T�i���D.=����M��b�4�ܳ�E�� ky��+��NB_S�/BB.�j6��_�'q܌ٚ9j��}W	�AcTq�S�:83�&��JBWO���@@E[]KkV.�1N�K&��>��ܚ<�Tm� 0�4S;jM�O�v��7�j&��,�pJ��Ooo�L�V�%Ϊ�q�[���,$xU�	Ɣժ��3jG&�u���p�Az��fRWK���SlB����b���X�pw�~a��f�B͐� A}c܉o@j?C�a��5w6,�����U��uq|���6��;�ӂ%�f�)�'壟"
=�\���p0� 8�o�����"�l�w��/
(�7VW{s1`�I%�,��6>���������nt��W÷]Ĉ�`</)�6%0���9�=�&�t���QS�4#����_̯�ez�Mû�k�,�
~<��C
���13"icIL���!.�.>rgFR��UF=��Q�G�
�̓�ږ�cmi.��J�,��3x���O�ǝ"T8�E���1������7]:�0<`��9�7��f��!m�u�����u,�.zӰ?Gƒ�S�\����/W��it�<�nU{�@�T���I�^�~�\o��\������H_��щ�]Y�qN�fͥ�n��pG���j��OS�Ħ�_X����>M�OR��8�]�jj@�p�DiI�|P���@v.|�@B��9ɹVK��I�4�f��[���裯�.�Lk�� �	�2f�M06q��y����`&��pg��x6�鞢�����O��x�H���d�-�-��A%* �$9vd�M �p���I�F{���\\��bG�����-,3��ul+:7ύ0G��؁�Mn��{w��YC����w�Qs��(�������u.s�!7�0MS\���H����xK\h������f���Sn��p[�+�,�^�k6��ө���x�1������q� e�F�|���ֶ��.Bl�-�&S����9e��S���x��]�{:�Լ���N�Ѭ��2�U~ė�4�x�z�Tȟe�f�h�)�k�l�����K�D��ǋ�z�f�j�6�� f��]x2��	b��ӵn�fa b�)�"k���Hv!� ���"�u`>��i�/� o�Sĸ��6Z�i����t��
���s��{w�r�~EAț@율���)�H?ôp?��	.o7�Q6L���Cf	TJ���FrK�X	����ǋ��T��Ϟ�  (d�H��M'ʬl���Zf����_�� XD}���}�_�c&��\y��%��s^)������2�c��$�;�skH;�Ő ���Il��D4����]ML�ǕFl}�'�$�|s�c��/��8;��:0���9�X}A�aKG^Ӛ`~~�6Z�:[V��*+�k;�~/�{%�vϟi���Q��,t�\y;��׬0�f' �d�� �M���0��t�ǹ5�O� ��y
�u ��[*ǲғ���9�\�i�������*�U�Ԓkfo��K)x^�0��7_My|ج�̞x��5Ox�9Y�#��psd��ȭ�_��yN�F�ꄱ)�AѴ���(�_����,E��m�dT!�h�E����g{ng�Xz�����^����?���e��M���4���k ��i�O�y!�a46Q�2"����l��� >�Hr�4\��%Sj:>$��y��Nd�������#�q�$�]�%�@�1}������lh�Sy}hOb�UC�X����Wٝ�{�8+,:ǌ��N_Z�nfuy�1kz���V#S<{���2a�;��Q 8�>&�'��A]a+���k�G�y�aУ��~̇ݮ���|CQg(��F��|�H�$�����g�T<�Z�/E�VR"�r�+^�_����@���#8�ꛠ�#uTd�$�Eف�