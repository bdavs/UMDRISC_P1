XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����1TUQ%���N��I\�!��2���� vĈ���W��]�'l�A���w-�P������.-��¬��9��]D��,(��`��G+���M�s�1ܖ�c�k��������AX�~��L�3I�N�����L�NJ�8X�4s�p�l����UK�v�g�\�8��"�AYXYj���k�8AL$7��_8������1��	pm1,gv��X��X����-�u��Ղ����F�7O��b�5��"ba��o�C%|�h2_��П�|S�*6�A�n�caK�$�I��>w�)@j����B��f�G��ƘB��mV�ᶵ���`]�d���Ȉ�ӹ�>�9,�s�~��IC~4�ku�d?���e��>�����n]��������ב8����0Q�ԕ���HX�'�/�gh��2�+rQ*{�|�k�˽�`bތ7��*0 �"�Z��"�h�U'?8'���-�u]]���tWZ�!�!�UGaF���<[��d}�l��nR�Owmq�Z����M[ǬZ�C�)��r�����ֻ���t'�۰�0�Q-�P[�c��^C�k�Yj[�6PU���WE�#�Γz���#�Y����-'+�ۑ_���$א�'��S�ԑ��.�9�$�o��5N�{<�x$���\��$!�Н��[�2��G�'�v��01�z#ydIv���-���z�،�lnӻB����PAăW�m��`{���<��۔�%e�W2��ET���eC2x��yXlxVHYEB    ea93    1880�[{K�X+s���X���
��R�5�t,
��#X�ʒ������tL%G����7�a���FkQʑ������[��c��l>�X������v�\65 �f��,ao�g����T���[i]���9m�ν�e����@�ܶi�Q/��Y�Ix"~M���V��J4��,�yז�Q}��)�V� j��oTސ;v�8�I�j_?"�x��I62}��O��s8�#�ј�.��	�D�W�dži�)~D)��'����9Y;V��:vwU���Sz�3.��gE�"Og����#C;%�G��"ɕ=;����*}�ʥҐ᪒	�G�wgU?(��M��k����8�sZ�3�����4�X�1�gHU�pI�~i�9�[���d���z�y6i�m4�#�3����۝��]4��$?��nO��jY���"q���lf
��dv���5T�9d!Z8"�Jf��C��LG����y; n7�Җ~C�Ae���>Δ�TB�mM|��yj���j�l<�+_>oU�i�j�}�}��u*���_�m�. I+�ر3<�Cص�4RK�|X�P'UD����x�)܎�!~`B��WaI�^�m2;ĩe����wh�&��_Y!�`&i>�t�sס���it�Z���*m+ٜ��5�5G�i��fw"'��<���,��AsO2���ܯ��\�naM8��E��[t>��}��:��5RgH\�Ac~´�;��tSD5��{���=��Z*�|qM\z�fp���U.͉uKA6���dj����^�~���\E?���4��^�����k6\�/�>2.h��5I��K�U�";#����O�'��O��dA�*�9�^K׀�����3�9j�e�f�Uqu��;/t0j"<�������_OM�U�My�ӽ��&�|ߺjz�Mp"�2�k��S���4,#�C�d�ȥ����5�n]��m���6((��@��بz���4H�kbÝ��KM��u�T�>������I�mfv�/DM���\�ç���dI����y����n���wƉ�Z�	]0�Y ��b�8	�BE�٣Qj��M�U�S�#�:�<ρ���Os���IOJQ,�/ދ�h����@w�D�����̳ܪ��tC)eq��3~�[|c��%�v�P����sOi$8����A>�a���C�"nw��P���p�(�	�T�g���x����q;�S�ei7h Zh��6?U��o��wmӗ�����kq�wJ��Q��o��W�ξ���t�ׯF�I����1�[�LlCI�$�Cy���B@�qu����^�v|�"p ih[Z����{���JM��@��A�аSﵿ�Rp0��?8/*�
'�%�h������TL�@��Bj��-�:x�.0��2SH�|�&$��ۯG��y���<{0���&$r[�����8*$3t����p�J��
����G^:!�n�-�N�l�[��a5v��,�ޚ�V�f�[X��,��I���>�B�Fc��@sT�y��:��$q�s�9��� l���1N����C2�*7���J��2_A�6M� +�E��_��'�G���t��<UWd�v�f�d�"��`@eY�(S}k����^3Fw���V��m�V�>c�N�=��z�*(T�}��#�坺��O��������V���W�y�N��cf^���Wq#�����0T� ��*�׻J��l�X튲v
��V��[>kU�v�*f�E�i7����7�k5�eU9��G�G�u|��l�v�lu_ K{��	�>~���ˀn?w}	R�!S����O�䰦�nnY!�r��k�~%,�lE���*�ȫc�S��^�Q"��ǒc�Z>4�0�{j�=�����h 
Z��$�����~rZ#���u:�PƢ��Nxk�s��?��Ն����lU���&�+�v%��MH���������3�N�S��_�]K�[�i!>����NJ��b����H�	�����0��@џ���0uV��x��5-��I�Xމ]RQq%���Y,�sk���݂�.ġ��X͏= �W�����<��m���U&l�UR��_WK���p�Cۅ�*|����<w�Yw�] �2���M������-��ŁYB0�f?���3�0i{�wejJy��ڱ/�MF�s��)w��/�:���{1S�G(��\��L*�M����>s�
ʅ}��� e�y��,��,��4��*-�n��I� ���L` J�,ܩI��\J���='{W��W�Q�ܳ8������D{����eJP[܉���YG�S9��!*�I������5兩5�/5�_s\�;��E�Y�Mآ�}li�b����u]��sA<W�^��dRb�����n��T�<n�Md�8 ��}bY;����#�i+$	��\��ʓ����G&��-!���<�"�9��_��`�0Ft;���v�K��^aQ`.6���(�t�;�B����̒�C1X�܊STG��
���i�JD�������y�r��m���Sf�Sw��n3�:g-��:w)0���(p�n�a����$P��䋎�&���),��޻�i��0��)n4���1�w�H�/Ϣ���+�g�뫶�3��0о�u�Z2�7���}~��8�t�9��&�J��Y�<++r������1�E�	@�ۖ�Q����؛� É�(�nܡ��E�U�L�Ol��ֵ::Yaр$���%@}�Ѵ�����a�5����k�x�,Ϙ�ʙ�oI2}ܼ�n5iå��<m֭�tt���HY���J�v{�ۖ�땺���X$V*�p�-�L�&��St9�@��Z��P��4�3���J��zsU�s���JAM���[᱖��n���Βo郌�2��8�cS=3A;`�dwז�׼���Zz��i�dfk���$ߏ����UԻ���*>/����x){���o���e�'?�hT���e�"#���;4,�3�Đ��a�6�:�����1^|�.��d���ٷj���ɰف�q�Cʣ��cڶ<��w��X^O�䐊�rC:3��l`B��l��Ш��l��������&��Џ����������8��ҳ�궆���%�C!�o?��l
Ĺg/T+>��J�v��kᗨ;b:k��|��N�(�����H0~빆>�:5v�=E`{�|^eMʤiv��#:��+@�
��D�ioO����2#�(Q�S���{�������z�P$r�ltc�����T�_�n�<��_D��k�<�O%T1���@]ܷ�^�n�m:����P��ڏ�s�����;��Ij)�~%�~Β��,;�Q&�mK�|ۚo��
�G���Ȏj�:���KS��	�z*$y�������cE0Q�?�[_�sL��[��G#�U��Z��%���ױ�^�c���1�=���J��ǰgd0����`��1H���4�����GA�՚��ia��'��DL���F�w� B�^65N��ҡX�ɱ�9��������
��$��<����s��_��cK�EZ<�FO�ֹg�R{I��,�eq��L����4�ƙ��K��[���ί����j���ȋe�45GRB!�y�tM�5�uM��R�l�)*�ϗ�I��IUiρ��K�5��(�E��W�[��+���;�D+�+��_���a�yNi|=I	k��-W�BmWEN��i�'two��W�rg��-+tM/H\��dr�oفs��X�u7�X����(�V:g�ګi�ޢ�1�{��J}�� �t�0��Ͳ�em�}�Y]�&������5��͜C��:}7�wb� ��Uխ���	�5'g�dv��NΆ]/�F��w��{J������(q��C��!%��Ξ�ܑ�L�pyTWy��5C�@���H�'3�V�O���Ș�\�E3��g�>�������'X-���ŉ
�u`�S�hߨ���Eӊ<�h��Z����n�\�*A�R�"�{c�1�z�׽��v��<�+��?
9��7ԟ`0 +_l(5ߢi����O�<��h&��|z�F毎��;�E���(�q���9-ټ~�Ԁ����@jo?f{�30
n�Y� �AS&����L�w�0ҭ���]���-�I�t a�`x?=�Nv� |R�}b�D�������1ϒ�eC�������b��B�~~A0�M���9 t�Oޱ��{J[�V�$�L(Q`�OL�9=�RP�})�x�¶�g^a��%�U��䟎�Fx���0�v����)���v�,{��Ha�@|�$��d�g�Ady0��T��/!�k�������'�W(�-�\�l�ؠ�����᝖_T��,���`��XA^��o���ʻ�^0�Y�% m�P'`��Ӓ���G�!�u�2\o3�3�0N:����ܒ�N�o��3�IH$]�R�+�Ҫ# �D��֜�8ؿ���(�za+�b�u�2ۡ��{�#f��a����|�K��J�&��D���G�����e�ސ���A`�N�UT�'�hp�u�Q�Wu�E�_5fR^5#�2jNL�)�pi�3�K,{Ωin(�z�qK���S4C�Gff�sV)9T�:L�ƇzE�wtӹ��F�v*�^�;�.^[�w����r�����X�V�&��s���s���ߠ��? �b�?N��A�i�t��X�	H��m(;Zz���+�Y.V��XJ��չ���ȍ� �ɉ�zf}�Y�ؒ����T�z4U�4m�z�gF\(X�6�#4ʼ�.
x4�WM,�Ub�"ͤ킷f��_����f��H���_=P&���P3���琹�_T4HK�
�Z���e���Ͷ���#4#�x,�t��[f�w�)��ؓ$gFL8T�0|,�t9��E�����2Ik<.�G���Q�ϞrT�a`�	>���n%��7�_�8�E����������+�r�ܣilP���D��Z�j4�P0@��3��y�~#��Vv/���C�r����ZQ̃- L �ؿ�
����L��h�T1��sz��&�����P��/�i#62�;*�l¾n��U�!���^<\L�%m¶]CM�ﰾQ�p?i�-���
����'|k3�8��p��H���Wtރ��s�!`�ֆ�����/��;M���DJ���?�mǁ���6�)��6�ՙ��$sQb�m��f�^�8��2,�R$ݯ�:V|�����Ձ#����"�����*ĄBN�_��R8R%kE4�R�?�{f�92�3l2�Y��YC�j�jքa�	3+,��Ǩ�3.`�O˺��4�B���ԯ.�Lӫ���ն�#;��2+˚��L1�14'�\ ��[��O�Ψe_qaaI51(�̿n��°3����s(�������MY�S%.�/���H�"��������7I��l�Ǩ1��O���g��T#4�ߺ?�NE����R��I�����M�Pv���%�����r�Cg�jǝYy��&��O�N��ލ�"��6��y|��;�#Uz�\6	ųU�U't;*�ܿ�x@�c�;�r��Sͽ��U�hDLɳ�Zfl~��]CO`�zzf	�T�R^!�5׼�C6�A�lR>v�;oL�o���;��R���Zj?i�e��n�߲	T <�#��;F)��u��E}�VM*��rd\�R�)�&�R>�[�N���Vͪ��`x>�:�d�5	�]�'��m�1� \��ke�'`\K����'c�Vn�]:*1�i�A�Ҽ[�fqY� a̚Ȅ2�%q���,������ٚ���v9�k$�"9��.��۳����$�(��#�ݲI5KE:A$����Kcciw�eUE�uq;��C�qf"?m`e�.>m}���������@�l-�BS[VBOg�`}���*<�J�N�6�q�ctf�h�e i�Q@�ۛ~�G�j�9�I@V_��+����ig�G����\��	&v�拱F*�Ǐ�;�G(��|cM�kQ���кR�	��^�u�ͦ
	�����A�e�?�1&��$���ˤp'��7�����h�FY����z�3�܇F�Mb6f�1>_��r�#?��&��:���<m+���ώ�kr��n�-zF����[��6p|:�WB�ϯR�?0��Zs�s���3�h:��2ir�2��돓`��