XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0��@/	��4'�.���8���{v���K���"��b,i���("	p#�U��!͆�)a'|��|��T+)a�!��s���"�����҄�Wv��p��a��j	Sh�$����y�M8� j�qS����l�� ���CX��}��ﰳ��SǬ�m'EK^��>T��G�|�f���4T�^����4<��S ,���#M_�&��l%��g=���Vz����R
��;�2A���Al\���+��uU:�E��$Lg)s�օ@���N���*J`XRH�աs<�7�"վW8/�"����}W� �ˡL�Kw��V��Q�#h�`}�ץ�����d}��K�rpR��.�kU��'ݺ�Y��E{)�	��/E|`3�Ĭ\���r���0��1g�i9~Ҹ����=Q�Cy1���6T�L+��ޓ�
/z�B]Z��/D>{Giz>�<J�&e��5���ȩ���R�����BE�E�D?Q+	�=�\"ZJ}c�e��MK�q\�Z7��q��RM����G��kϥSLB�|A{�B�@K��7����=��c0�Z�GW�s`͢K���E�g�o��Y�^4r+E������-�i׿�Ԃ��-ϴ.|��1��B�����E�8(�<���.ź��i��@��=�Gq2������se��Z��io�$�5�1�Ϸrq7}��|Q��9��u���B����_�[�Z
<v�6��l��൧S��XlxVHYEB    2e55     b00��Ձf��z��̂���`�KҼ>)�<*W�i�j�^�o}5�e���m�V6�����DDi�0���+��M,�3�sy�6Jcb�����:�s�)���6��y��J�`���g��gH���ث]���X�`$˰�&`�2�q�?�"IRL}����j&��k�Z���dsv)��#��ݗ����2�?0;�j������K��FA^�C��k�4�y,�"ut=￫�O���I�9Q�b��R�f��T�k�H&�5$�e3��:��'{��9�mw�r�?p|2��^	DS֠� ���R˷A�5��?r��0������v�R��yI�����"5��A;|*N-khr�fs|�ov>�L���hH��r56o�������*�qҬ���ZG�a�%ƫ&�NU��E�	pGy:*��RB�7�Am-��bc5^X�H�e�ͪ;�$?_�����xǤg�7,�K^"N��N �ܛ+Kw�v�N��,`wv�BWQ84[����Tjh�����P�M��Y��N�.������`ҷ��O�1�!�9w'��z���ʠ���W�#�:�'�W����|��@t/�+utm������}�. + 3o�in����t���0��F�8��7Ukdl����>^�:>w��h4�w��8��Cj���X���|eJ�h*�7���S��
҈�{�U���~��θ�&;H%�8�����x�Xh�7G����GcI�p��>pk�����l�Cُ��}�d�`ҍ��[��r|Q�v�3Q���3E�X�[�	�Mg߲�pF��LM�P �R�X����2�}|lS��٨U�<-\S9]/�`%���Z�A�K�ұ�|Q�э��Uoru.W��T�q�9��~E ����V��2PqB�PO$:62��PM�����}-��)�Qn{G �DF)�����\��X�F�{sErr=pliZ����C7�.,&�$�
���ز$i8[U�X:Df�rZ
_|��
\��;�U�r]K'Q9�3.�`J;�N�9��7N��-|�>��x!c�,��)ݍ����ޟ<��q!���@�pe��C�l�����{���7��*V�ɸ��_k�-����w*?�K��WS��0F��7�&6 ��yc�</t�hy��q�КPR������t�(�#{��3.3��Q�B�P}~�߷�Rv��~�fq�;�3Q�I��E���~�g�S��~�d"'�qR���%6s��&��PADI&��,�d��a�AV؇Ѥg�z.f}#:7�K#��kҌ���.5���5��0k���!툏ĖO|�p���p7�{�tbh�-F)��\�w\A�WH6��P�ئOe(�E+�.X�tQ#'P�
�!�5b��
�$�B�c]8��Bb5�PF�
��L�F�}��l�F#t��.�H
� ����2h�ħ#��c�U�Wr�/��J�^��DY��j���I��' �{�ꘃ����$���E�%����*�h�� ����G|+ly|��c��ڟ�_�-�����M!Cv����@\��2�Os��>�B`@Sy\�	FQo�w�mE�<�VpD��O�Fvg�@�s�۾�;�!��o��O�i�N�5X�0�}.�:�W� �:	:x�/���E=�@�D�8ӫ���rO����T�X0�;Eg.�[!`�4�����U��W��3�j�r� �p�d�B9��;Ҹ�OE �V$An�X�.���(����g$�P��:6F$�@�ځ�Ф,P��2MS_��l�4�V�808:'�[�5�ȩA)���6F�G
���4 �8���w�]�&�Q�%S|,�|MN#��5��hɍ[��h�m`�3�}'�Bw��YA�E^V�,�����Ҩw���D͆b�t¹��GC�m�5&n�n��@���dBA�k!��^��٤(�L�X�'�!��!cJYt��<1,�2ʹ�0��mƄT_���bnR�d�Њx� �����y���[Ѝ�<%�ͺya��]�(k��R�F���%�g�q^㍶4�����,��M!"稐b�r���``��/�=%��;��ڄ,�?�D�痜�;)L�_T����yY �iy{�TWJ	�\�DJ25e.e��@k�C2����� (�_�%F�k�\������ypZ�`(��]j��.�c�%�)"�=E�U]f� �s��8}�Nk��VCy����8�������{Mvz��2����"��������:���_|e,h��%�H�$ ��v&yT�}���%6Z�.�Q�#��R(䆳��Ϗ���Ӽ�(�d�À�U�\*0��x���N��F�E6�-�gJ�uV���������].�ю�g�RgL�m�!��|O6���1��4"!U#�=c�X�\�"��w
oS^����������㏆�GI���Z�z-n��d��W�G���y��{��|/c��1����0�V�T�'B�惨��0*����&�@�����Ope�7��>v�9�c�4��-�\l�0e�=��Q���l$Te�M�W4.B�[�&zMst3ii����?���obSp�2�ߜ�ٸR�D�7|x�_�fMR,F��ܡ���s;�� U؍�F��8Jo�|�)
G��ݸ1��Q���v�n@���X�_8��p�Za�R�!�̝��+H'K`�;n^�N7�Z=i�:�" �mn�����Cz��g�S:G�ǲɵ`bO���b��z �[�W���pgR�)�O�n�m���E��������1���+�i�Mi{�	{xƮ�V���_���[�4�sx~s��)�[���O