XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W��i3�]D�U��\�}��N3	3*�����������Np�%!F��p�6��/�W��O���!**|z��������s�| �e���=�4 ��he�N��M�s�6�f?s9��%}Ӷ0�!T�tTA!�d�iX���Ĥ$u�͛47�h�N�����/_3�;��]�{���K�����L�"�Z��GaZ	�4C"�4��pr���a����3��Cğ@"�Qk#�7������+0��uW�>
L&���'��K��>u��{��%v��*<�<J�8���]�؃M�������9�h�T��Z_�T�<0 ��-�o���I�Q�h���^u��=�y���MɆ�nٜ�Ѻ�&��QU��dY�jvfjm��M�I�M|���y[��s^��_ś^�"��>�L�!��8�y�,'���G�}]�1����v��2�~���c�z��'q�A�x7��C���>�C9�̆3ش�M;� @ɭ��ƜGtf,_�������Q��Y��S>��G�J�D������@4%Q�􂑰.e�'z]��DTNR�("U�#��+m���n���@B����F7o�[� �(u����!:s҃]�����y
	��?���!��̏Y7����O�C�.b�#��4Ե+G��jk~�	�4�\d㲓��D5��%�uw������@���J�kݞT���y�']��P9]���Ok-|rw�>�s�X��V��=������b�D�T /��+�%嶠�XlxVHYEB    fa00    2480tNߖP]?`n��>f���VZxF�Iܕ:[�]HRs�[c�]j��Τ�<�6'��i\ϭ�V��^$���l~�;����sq��ũ�1���+z�F�~�a9�L7����+%*X�"�:{95\�\�鋤��F�D4nC?��~�I��E�
X]nc���f.���4�0YC�$��0�m��Kgj3��@��7��n%��g�U�� 9�֦���w��1s��R(ܘ+;3���$�,�����啌a{\��Yqi�B�Hߛ^�(��]�:�4��Tl�m��zA�*�c0
����H�1$�.�V�+>e�E3f7օ1W��T8���Ӑ�Y�p�PO�j�s�}}0�BN����k'�������4$+�����%y���L�t��̎���i�#P��}�3�P���÷b�oϻ���� )gp�s��SF!�A�1���CQ��t���]���AB�$�Mx_sK�:�e�^p	J��A9��k
�k�^U�$�N��y�vA9��ʰ�dbۀ������3K�u��\��zY`�$�E��:���9��%��d~�Ŀ
7���x���0����Oe�M�͢��^���)�sQ���=r�y���H�'|!|8�t^�_��*y�� ��6�3��i �Rў=Һ��6ñ�DqV�r����U}���'�"�ƿ�0��w�jG���]��i�k<���|��K��-Z��h5\^k�)����*��cu'v��(/ �����˫�#�y}u%��;������3#�T�u����t��	]t�q�p�_��'��P���>�؆�4T��֝�@~���e�~�n��3���`3[�I�Pw裇V��u�����"��$C�S����]�)��j�Y��"qÁ}~�����C�
#�t�����;�蝹N�vy�Wh�^
�@�V��0zb�x#I�)�!nƼ�xÎ0�3� x*��4e���Dd��Pr3��o���]5A��v�dZY����	^�5(���([:f(���[����[b�M�!r��T�ڷ��;Y-�J���,6���/�=|̂���E�~qgR����}PI4FZe�Z����d9��ϣd�7X���U@��v�R��_�&�}��=DH{yl����@�?��!��p0��km�0�����O���E#��6Ԕ()�����d����4�� 6�Tί-v�~$Dz�l�ח���0[D��fޝ���.�ؐ���M^�(G\�!�i�[#��/����D�����ѐ�T�N1AZ������{�ݟ"�Ee(�!���r%~okM�)
��G�6G��
0��G���� ��h]�g����5����aP����e���
�"�	[����eg��DA ��g�I`��k�j�%�+���ʹ�P��9�g��F ��Ϟ�IV�a�$&pLsvG�(��_~(%�0e�����=�/7Bz��J	.�[i��"&�GD�I��s-CL�+4(��Zqc*X�CG�>�ŢU�y*�Ȉ]��5�^O��`�԰8'P�!��(����(��f���,����N�1���;��fF\+-�2�o�{[��`�l���d�H��%���0`�����O���l�2x�����k�j�ݸu���Y��b��߬,�NʴyY �:[{Yp���ay�k0��#-��'vĹ����0FY�}��K��ꇦ� �O��ek�f�0�Vm�9�h��Ӑ?�n����<L��XEk��8X�~�����\�*��3CJн�7�r�	ʨ��^��	4����`=�0�]��c�A��tp��Z2}�p��J�I8�H���QR�c�8�~f&wۖ��E�~�ahKB$���ȗUh���D!��� ������<q"��q������~���r*vzh�n ;��bx"�4<�I�G��!�+��@��ˍ�3
5\��s� m���zuW)ߋo�_��a,l�i�m���,���Eԝ^Q�h�ܶnڭ�8>�d�w?����%��N��.�x��c�kb�=�����Y�R���a/���Ma���:��,�aY��<b����]%��48�kb!�O���i��}P/'t�b����,l+�RL�0��D#��k�գ�B@?�%&>n�B��s�a��
�E/��FP������:.��1�h�R�{�a)9b���ۆ�U@�s�3_z���%?�J��J�4��4\�ht���Bs4E��1���Z�1�Q%��<�#�����%㛾x=��e�k��y7%���A�J�J����j򪣁���&�êu,�½�w�D>�.��(�� %��ѕr���5J�e�Ɯ�{r���3� 9������CCM�m<��&�`�&KV���ĺas�tP_e�)��H�3�َ.\ DU K.��5�M�����u�́B���Ǽq�/(�̕��1_QЖ]Ue岿n�� Ճ�yB
t���3��|�׼<a���GZ]p�^сqM�"�+ٵE{9K�b	�5&M�oK}�I��đ-�K����eY�!��d 	�
�T��C(��]���|iIE����4ݹY_�	�=��$E>���BdH�����t�: ]i�_`֌��np���q���^�����[�g��>OfUw�#t��Ef��'b����x�jE�S&��D�Vs�6�$j� �9����(nY�Q�u���юӔ�6c1�Ŧ}fp[A81�z�ލ�\' Ti�T���F�(��j,�|���J*�i��G$=�[�PC�,�8,X��r�%v��3��Nc���U瀙84�eρ$ӪqL�mj�h�UVW�0@_�<|��א���w��fx�#hg�ڵ��X����@���v�^Y{�~��+�H<뼵���g����T�Hp��4����3cE7�PB��a}�n+��18�_��������ӝ��>�כn���ӻb��M������,�����tfu��%�M�{#��v��V?���(Z���5��J�����
,��LPκ�p��P�}���*LQ�@Qg��]����&�"��B|��dQ:|8
�x��uzph�Ň�����k���:�bF��N���Ѽ\Vf��:z����Y��x��	7�b�\;��T���.�!�v�ʹQ�交���7�w�l��S�I����'�����	4h}g�v�үy�����d#O�A����F)*É�w愬�
i�L�
R�6o�Y��'꯼�©�镣��gI@�q���3-�zF؄���d��V�j��|&k���τj	��X�Z&����s7G&GR5��mF9�Լx����*�`�Ǔ)iwT��=��͕�ڥ�?�,"�-=$����Q9#�ƀ��XC��F�y�0d:���F���{cf�Q}S'o"ǜ��y����� ZK\�|#���"Bs����ڰ�G!�XϦn9T僑�"Ȍ�1���:�#vg���PR�Cs���	��=N���P
�۴Q�g����V��Ϫ����n2�5W� !�u��M�i�I�6ʄ�{��eOr����Ј~�w��Q	�El�����)�]���j�Dd�:�%����|H'BJU��:w0����x�.�N#G��^�ޏA�H����:f{[�Y������ҭh޲rh���k�[��.ڴw"T�ב���v��`������U*�!�e�(�fZ�g��M���K�	�u����q:L4ǾS-$;,�f/��l~~7���
�_yK�O�ē�LV_SC�kϫ��NzP/w�Pq�{�]u�."���z�W:�;Nzj��>�� �9�h�N�H5u]���/>Ph x��>��r��tc�K|���`����k�i8�dD7�8�B�5��4��
'0=��Ǚ]",����"�%���+����P�b�gޠ�P�ؼ�-A>����k�������:�;Ѵ��������5�3A���������`�a>%�W�"�2t�N�<.�MU;���������ѓ�����vF��z��(��^:
�Np�|��3����y��y۴G{�7�_v�`琱�_\�M����30y?�X48)g�/La�>��	$�@�Y�8��#�����''��Z�h�7ˡZn�/��:n����N'�?���t9����&H���>yM�?_/��j�V����9����)E��}�ͻ�rv�y�u�𣿋�*#xȜE�5#��+3*�o`��D�ܞ�C�w"�>[l��[�O��
gz1���F|L�ir�~��Wz|Y�L�b�?"�l���f�xO>%����hr�~"�Z�&g��H� ��ؗ��n d�[<0	$,�9ԆA�=X�,Y��~8?�<*�mcD��-�*Z�&�W�=��wZ�{�r�;��`ʓ�7��8�;���Jf� �
�FȒ����F	{�w��l��&%���Xe��N�ꥑ�V������*gǼ�fI>i�Ca��V-���Vh1��vi!��?���J�.F0��SJ2���{�8�p��),��%�9y���O6
�`_�ԅ#Q�{�g�9�0-4�S�P�;ϝ���{!֐�Z��|��]�9��p��5�r���y��R�)���Os�cvO<�xP����AQ�<�ɨYY�+����I��@�����b�阬��P���1ok���к����P������V>Պ�v����X1O��2�Z�Vy�7
�<A �$���(�U����"���5����d�g	���X��!��J��*Riz�i;kfD`5�bZAex���׫�CK��L�L�Q�F
F�!�
�����{2W��'�8� X@�,��b與�d�����(/P1֓���v&@F做�*���_HI�;A�u'W<-�Pm�	-��l�P�e'W�b7�b����A��Y� �9���)��A{��N|���\���hMc��B
̤&6�bR(��o۱��)-���W�Lx�b�m��>���Y���!�k[�!���6��3�Nfޒ������v|ՆZ.��iJ����W���I���"��,qv�� �p�p@�@%1���J�N�w��e�d5+/A��3[�T��(���,���#�gv?�9z��7S*
⎸9A}�Kq�Z*���� I��Ϲ!	6��t���"���i�����T�>�XÚ랹�����Cg�m<N�gw�i��S��켩���b���s~���#�89���0RÇ���@(&�'WI��ګ�	M�c�_)#�<F�)�h�K���e�"������N�"3���O�^��=�58�D�1�狧�&�9�rGԷkC�!��BO���}c�A��ԁQ{���glڲ1�Mb)����������6:��aJ}����s[�5�3^���bnl��q,}��.���9�,���b.M����ĳ�A���8{V�%�VÜj0�xZ̖��M��i�%��G�x�n�H.��+�:{�Y<Ʀ����4#�w�x�r�뿻�s+�G'�	6ǿI�����j;$�: �E�v͞j}�̃�[q�[م�f��~��>���GU���/\9�UpNfh��Y$����5�̘�Ȁ�aC��mO�l��si��M1)��.�!e�Sj5�=Z�WB�SN�00�+�(����GO̹�aX�	�N����@�2�Ꮭ���JV��nMW|D砘G^q��d�X(��^�U�&&�zNV��/M��q��i���h�W������9�5�����4t�ī⦲��������\Q2^,X�������6��qZ��$Oլ�o����F@$q�{�hva��}M�UX53H^�(�K�A����A��~Dl>6��J9��h��Ǉ���v�;\Y�c<��B�����2��f������t�r�=ڌ�ȣ�O���Aar��"��L��5�I����ޚ����vB�k�4I��:��/� ��V���y�c��ݠ���$���;ǣ2���o����MP&i�W��z��a�~m��Y�[A�G��RKޖ&�ǃD�� ���D�'�D򕛩�=�����kܢkL~@QU�.s0�={A_w@rv@+�N�.px�sޡ�g���^��j����Ё�h��3`��'���s*+&�?Y��7n���d��Zؙ6�����iZ��z��~3�#Mx���y�K�5I�%�A}��6U8U��a-�6���8'�����{;?�1	�)t��@����qd�q82S��6����>��qT����T}��'N���uG!�t~]�< �f����Y�Gp_�S�̆��D�7����-�ߗEp�u����l�mJ��ɰ�w��o<h�wgx$.����W��n%�Z(�@En��A�S�������K�E�O�.n$��O\y��_�n:�nL�G�`���
82�8dUCg@�o��d�P�����f�D�5�5���*����n"n����(D�0�(��� �	��	�\R�n	V����dG�촘F��&���=E��a���`-���'��ۤ�*�B5��֔e��Q8��%�_ �ٻu<�I%�/�ʖT	e:�T����V��Ԗz~�B�M>��{֟���L`b�h��O%����,�\��N~���R��1����o21���{�7��XH6�ᎇ��=�ρ��Y7,�VzpF��-R�][�;Ⱦ���LʄލZi��sGl��
d9h��9�uή�\�jF7>��E{��=�U��(�Bw����2c'ښx��� g��*����B��A���X
>p�y��JD��5�o�,���ZpB"��S$;c�-ij�e���5�
����rIr"���X�����O͸����W����O>�vc6ߪ>�B�J@;���I�]�[�Yi����;#i��p�l��W}���U�]��I0s�J��~�!(/M$Q���RMs�y�V��� ����][�N[�ހ[���C>������S�8Ij��9������~� ~�oyD0��^���x0D6mψ}FKyo}��l��K�r�P�e*��\
�p*�7��O5�<�O\
��-R���x)�I��/��P{��b�|h+T�֮P����/K�=_bg sv�fG9�WS�Z�!�7đ:���Zi�5>c+�,3��j��2R�V/��J�z��4(S(�Py��v(�+�Al��xr��`5�va
���i/��Q��~����zp\�_�4���n/�es�E410h�c(�7��k�;�/(ugpa�Qj4$@($<�13'�ʲ�!��i�Z����H������|�ǡ3	��c!��ȞT��}չ��V?�ޮS"�|#	��o��Ư�Ķ�V�\�_4P�r����:�UΤj�L6A~z����Nr2[������d���^����ܦcIb�"���R���d5f�a�a�ml�����pb1�"D����4���-)�kB3�,�q'��ߋl��6�x�����yU�=Y�a������I�\v��jP���ը��&Y�vȫ/���sj��a��M�׃��F+��+T#%��Ǹ����0ن�u��K�FP�g^�2WI,iLT�Ѯ\Y����rQ�%�y��F�7��{����ES� �`<)Ͽ�|�8���st�w?��m��vM�AA���Ӎ,� �6l/���xT�`�ĄRܦ�+�=��J�ց^3�K�o�%�%�R�tŅ+�԰���r�g�5R�����x��c�S������؀��|vM�)u`�$����}�����W[�CK�J�_'~XnW ~� `<,��6�-^�j��ώ�P��=iu��� ��X��d�i�yW�Bڔ2�]]LG^�5�s�n�w�DN�ɯ�E0p}3�K�>����qj����;V��/��D3���vL�b�6��Ԓ?ڮQ�#�+�0�����w���E�_�@�N�xc>ᰚ�������\���F2��u���r5t-�!�r�Y�7��.Ŧxo������}�[�2Q�.�Va�	Q#�Ի�H�J� NW/	�8 �sT�D6rf���Ϳ�5�ޏ���D�&3X{����2=����y�D]N���"!]&sI��[�X��fLH]��|Dk���R�P���xIt�R80a^��)��U%#hh6Uø��鑣0a-�0�d�]-KWj��ӗ�#}�D4���cA�+�*/9�T���O���Za�*�k�����^b8��H�AuXb��r��$�r Qu���}�g�)����%ٻ9|�M,�*|�5c� �9x������n�Ϣ&fru���
2���W��J~��b*��<&횡��,m�aK�@V�`i����귲!�1HD_� �:`Et���L,��q�PP��/��x<����fodBeē��+Ux��Y_'T���wQ��fz�T�j�����,�"��Vl��Fa�hX|��Ko��4�C�mGBkvm%Ɯ�G�9~�l��yC��
6o��Yoj?�%�f�!���́����P@	&Rg���$E7K��]��7>iB���c�<y�qE����@\�N�ζ�&*��O�VK{M[J��/���j���uh� ���L�F)<��]`��Nbm��Ҟm�q��	b���È�sh��8��E7�-N�y��A�}�o�R�v|�i��8��ˣG�"X����ڝz�id�߯K*M�m�+�3#��o����$�+�
��_�C�f��QB� m��b@
��N&~�=E�Ɲ��̛B-6Y�$�*Z=�����X!y��r�Lj��GW��j5�����F��C*��8	\0�Bi,��*�?=��Y�"֡�ꏞׄ�hxb��22��SXk���W f.�s����)7/�}��qr+�i��W�-�`LI��)+m��M�}X	ݡAK\���r��	Ӽ2�?ڊ[�L�Me�N��uB�ԑ2� ��̭������>���X��Èl��e���ϪX��lrs(��Fo��k��L�pF���Ɇz����,��株�Y���˝��/��!�e�M��j܇�Q_VE_���yԳ�����M�Կ��7�wǺ��#Q����'�$y��j���IG�2�z]c�8`�!��swplk�T���w�7B;%.&�Z	jU�,+S�����Tk'*����V�D���۔'��eQo��Ύ��3-���o�%�d���˓M����(�]�'�A�Q|�V����:�9�)�I��hK���	�S�l�|W�q������k)X�ۄe+����,<�XlxVHYEB    964e    1150�!�ۥ��Y�FL1����G�+s=o ���6�^>�>hk���Su�<k���1q��ʩi�6�|>I���i�ǻ`^�xS��n����
�X+,B���O0Ų���<��Jdo��p��� W�΢E[k�"�ȿ[ȅ�k��|���Z�nqM��1H3hTvk����R�ne�ٍW�� �L<��zU.<��>�3$�vD��k���+�p�-�HR(��h��/��%�B4�ݼ�u��)��Z�`+�o�n�pf6�|�����k�Q��>,��Q�
�B�P�H�_���&Q�j��iO�����r\��"^���غh����x6���u���`Զ���G��N���3����w��^qT6�]�;�@�\o�8���y��^�Ԓ
����ñ5�aW�x��
Hv�:���״iX�E�ʁ��UڲJ0��Z5LDW�١T�&j�S��d��u�O�y��WZ��cD���:ä�X���`���h��_�UC��($������IT��sDN��HȌ���"�t����XQa�"2s7�+��#� MU\/�/Jw��kr��;���Mzx�����^�%A�@[�ٚf:�>v�r�����n�-�}�~l��d������gց����`���w�X��_��_D�n{>Eݟ�m�g�em�Ȟ��u�ru�iF.��مZ��=j�p�I!��e݋�(t�)����=���,rC5,������E����Zb}����j�(��K�F�l�9��wR�!���CR/Z�Fn��� �[�d.�=�[@��O<Ǖ�r�lO0V�8��,�7���+�]I�9��12���8���.�Đ�c����
�x��?�J���U*��Kz�*c�ן�����V$����Jm�a2]���N�����J�1Y1���]mSM`"*�*=�4�V5�=��xZ�������C+�Y��f��\[{b���t���@�h	hb�O�ll#8���<4h�Aδ��I�=�h�G�`����1�ѥ�%�rd�*���h����t�,��m�0_Dk4;�w.[l'�e-�"�hK!��'��p�^܎��&0�AVf�:4���ѽ��0m�����Opb�1���>��"��o��Ѐo��%���FS)HJ�����K�6|m��e��k�!�f�yD4;<o@+��c���p�u�%��16I�}A�~p<h��Ɖ�g�9�EQ� �Wq���ȕ�4*)�ɺ�~�;������Z��6� x�w�h��˓Ѕ��](�=�Ʈ�ulwMW'k����aZ˭J�^����u�zU8���n�%�w�G��mǽSUQ���7�%#���;���	��Ԡi�~R��zp���T�dܣ@m���?'4M�pD�s�rup���m΂��!,�8[��G "��=�@�f������\`T�#ύ�9�w��i�,=@ز{
�q�`�F��l�����r�%�}a|���'�q�͕L�{oKǨ7ھg��ټ��)&���l�I�ZF]&K������vwV���DUV���r�#j��Q��Ʉ,L쒅�3��=`4g�(l�G��O����j�xj����7�i>���oY�ϿS�:��2�8�%�����u�1���@��j7Ǘn�Q:�r�Ě���g� ��T��ܪ��l�_9��ˌ�gP:0���:z`�;��\>�F��Y��&��iِ=��U��I0:���t��Pc�9s�⁧ȽF�~�<n�틬�t���)���\VP�ߖ����^�SN5��4
3�r��@�)���v����Ώ>�	P�%�{\U�`#��9�ļ\CDC�N`B:�K�Fb�Υ�-2h썮
}�e�)����W��q���\���b'��+�[�I?��pϕ�H�F�����h,�f>�kt���é
�\��/�T\&#�u�>����� [9�'M��Yrn�󀰫04F+�j��9&��V$�)�m���� �5�&4ı��~��1�-��o�\ꈳ�����.?�׶�����#	��ٵ�@ɐT������Lh��t9��_���_�
��f!�IHe!�����K�ڽa��v�$��^������R>&�lW���� ��->t^���-I�ZWճ��ȝq���Fpj��=��|��\�'��"=�T�궵7��������34G�vL�F"��ca�Ϩ�1�5Ɨ{���y�.ps�@8��~�bѻ�W�օڊ¼r���o��;en��ʹ�H�GT����?���|z\9��~Mx��wWX��6X���,578�ʛ� -G�lˢ6{�	��1��D���d�b=��y��}��O<�\�w$Sѣ�w� �z	��q����^ߴF��(�>�T�_	����~/o-{u�i�.����D_ʥe���ss��ip�Q��pe�4�2�&�75�$%����Z�0��k5��L?��dM��4 ��>pLn��9�BN�E��O y�쨉�_c���������7u*BjY��4A��e���2�y@�eq3��P��;���h�tэmz��K�i��(2��
�U�pM6a����EE0���j����m��:Ǜ���\���B��NS/`��S�y�C,$/��_Lg�]���\�K�hR8��6o&�_%Ƞ{ �+�fq��fW��7�����oɬfK�@����a��y��*�i�8R����������̯������g�P��	q��T����@�͒�W�h���|�3hw��e�*?�Y׽zO�\�"��ęx�U�[�-�ʱ�gߑZ��
��7\��ה���5_O�,���|*5j�T��ݷ�L�
=�!ǭ��;��п�T�UxJ��a��K�٭��.��˹�O`�]��c�*���OLCތ���*,W�r��۪fMS_U$ 'o�S�#ƷFl�C�ي �����]\f��%�����<h�f��*��
*�{B����킹��{q�_Yz���?�ԟ'�+�k����Q��U�\D���'��(a�7�J�%2���`�N9��|e��"+[#6����e�6՜�\^�OU)��u�#�X���f��|mJ8j�6��-x�P�@;v\I|2�'S�A�A ���2Bo�|L�*jz:߭'�9�hwD�f�u�Yy�(ֆ����B�����&��q�@�H���<�ށ��y0�?��ST[�_��D�M�u��m���_�r���Զ$jC,%	��5�%E��}�Jv����J�������RX��Ρ���~�݈����%8���D���o��h�2��w�G��|vZ5|W(@��Q8��tSo"X�=�����
�n<x��AԮ��Ԓv�{|���\�̘��m��*L|])ո��ȯv1�r�����6�r��s�/xJ�}+8�f�ӈ��k �\9���S�\j�n�OB]�w!b�=������V����]�E6��^<Q�&�@��f�����uͮ�m}{�~Bl��,��݉#<y")�y۱�)b�w��R2��.��	�����S�,�������]w���AC[q�r:���S���_`����UA��v���?Q*��!>�`)u�5�Ϝ�����x��JZ���nb�� ���a}V���?hѳ�������?�"ú6����Ȩ`�X��>��򘭫u��<d�]uBb�x������"qM��t" �����\Gf� H��u��/;^#%U�gMl\>3iv��d���RB���D�1�ጿ� ��l���y*��p���A��b�8V��G%rm[�pLu��x͞r��\��k��0�a��x�/sx�H��W��N0��ȣr2m��=�+����ɧ)��u�9��A�|��	X$��p���>.�kǮ��)��#v���U)(�V����z�RO���UY���I�;��F�]~��t� .��s�X��Z\���ӹr��`TQP����\�s65m�'Qћ�Q9���9��G����`I��")7���X��mX���.=�ݿMt�G0�(u��=��@X-�̷0�-�]���EN}�2�NXe%}�gB��7�{�+e�,���	�`�j�ms����h+�_T�#n]J��-�v�5
�d�_s�!���.�I��}=w$����?�_�l_�YZS�y�hEf6�ȱ{�M�:�BZ'�w��6��#��6%��/�Y
��bU���Ĝ��ɉ*z��/P�z�/�(�J4��� ���jH��~%�e˛�<�q�i�[oS��P���� k&g�Sy�Q�1m[�p�����5MA�������H1��[%�1�J�
�!
��