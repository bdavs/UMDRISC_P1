XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��It,"�sTl���ml߫@�31V���N�Ӓ�t�S+$aI}<�(l�F_���vFv���8�N�h
��n�/��ᅰ��ݪ��n��^>߉��Q�P޻]xX P\�b_��b��ٕ���Vq��+��%��/���-q H�=ˮw���f�M}��K����J6�]5����>`���䫜힔��Ͽa��O���W��#eF�O}i�`CN��M�>@�+�Q;+�4���ގ���Z�ǟE�{م� '�J��� �f(� ������t�A�sj�U���n�b�Nٳ�n�堯�k�m�#�P�!Gu��Б���f�L���ص�2�Z?!j��+Q�&'�&2�1�u)W		މ?��h��Vz*"�䦀����Un�i+�LP��n��M��e�����O��L�AKA? rT;�x������/�bcTDH+n(���|��Fn+��1����*F/�)З�����2�����8'@���o��1�ζ�S� �'�O��K�W��Q27�1�ucN�U;e�b�Ȕ=�������[�E����!���B�].�!s���M�����
�fă��n��=fWɪ��^�/���2�΋�l�7'�Q�듨�<���Q4�la֝:�!k=BJ��k �Fo0������'NgDe�pږ?"�o	�a�o�:
<���W?@��Rk���ҳ	J���o��*��V��� ��;�:Z�'�q[W����Xꖌ]�\?^M	�
2��j��K_��o��Ma�XlxVHYEB    3504     cb0�I��$P��Zo��MD�9�̜[�$�G|�[�o�<�2X�uf�2�:,D���R	��Mt�1�	u�)|
¶�x��%0@�	�!���49�J�U�D���|XbL�/W�� �qPl C�p�|Ʉ`/�oqlFtw,��u4��(��gՌ:C�#�S^\�]��?�������X���~�`6�DȏR{9+�}Y>�wgs�C�z��!����v��a�?#�3�&�ֵ�L�/�'�4
h�����1x��Q!VȐsH��vV&r=0�sՆ�s���1]˜Ň`���*Omث4���=��\��b�Vq���pc�`��j��V��0�n�v�� �7plX�l����3�a@a����%�N ������?��hM/z�i�!�<P��4z������;�E'���g�sY���ڹ��K��;Y��*&Ѽ��;���"P	������pcl	��/%�k�z��_gų�
`��g�M�u�$�qq��k���� �5n\Zz�����E�?DkT�f��TI��/AHm|Ȭ�(�"�
�24'�)n��}�a-SnN��zNc��L9&��X�Y�=]�;�2���F"J��d�E�}�Oe&�|
��`��ד�A���₇mV�ɳ�KI�ZA|�j(�A���#�J���Q��0�X��U�O�^β�S�q��u�uR��Tr[�3�a��<��9���*bg�:�L�~
~r����?��+7��
�^1��\E :=��d���[�d��N�	ObG�+��+N4mT>�`�,o�m�����ud40�ٕx���O�?�1.�֕�5� Jڂ��	qD�r	������a� IA��ʳ8�([�Z}!�S@�T�F�?�R�胥a���[\B�����`K�+����q�u���ݎɠr�^8�"p>$, 
ޥ�w�:�ol���+_�s܊(��w�h���x������w�\Ʌ�����j3c��w6m����1��p荒�wɭ��H+��0[�m����&5�x��3f_��`	n��9;��Z �����C0c�����!�V����`�N2hr�1_8��F'��YҌ*Hѡ�L��nlDĴ����KH������ɽ��_�z�2��_>�[�G�a�'�Ŕ �F��f3 ҥf����9�>�-��j����e�ew���S�;	��Y���*���͜;x��9��+�m�)��Eׄn���K������b�щ�.l~p
�5�}�"SOa���1j+�s�dHp��P_Ť5��B�����b��<eB	B66U�b��@h{/|�w�����h��A)k
�6��a�Һ��e�X�w=�dY��ۑ% ��1ǼjΜߔ��&V��֧D�[!�83����)�PP�����5��
6T$�u>s��P�N��EU�pp���=��Z��HD:+>�!�<�`�貮�lrÑ�m�h�)��n�)��#��[�t�M���z*�u�5]�$�ÍJ���ۖ�!���\���n��)�#��|�VY<4"!���no���]��w�#T~�i	U��ED����í�!=�|��H<���B��ر�~��$���b�W}�;��ȯ$�D�,޹QF�k�-٤�}3����q�8�E�L��R��ӽ�o{;�ң�c[uU�֌�gv2-�`"`�ٔR�����B�RL���u|����M�R܉@�y\��d�|�|�W��~5b�%���`@�<sc/%���hX��}[e~����[�:��rT�o'���A)^dٺ_u�����#O�mvCU�\sr�9Eba�մ8!_=����:���e��M��^UK�4�
ܫ?>}�t�{c>�؈��0sU�²��&�k:�X4��^1r\?Q�]q�:��ܐf>�GWh�8e��2`I���n���i��.��+DfO
�S[w�n](��+�E��ǅ���)B܋��-&�����u���S����c�R�ĭӵ^l�TnQރ��#�TE�Y�������22�ת��w��R��H��z������֑�.���ߞ���l&yp4�����^�o-(�,?b@���dH(`G�\�9l7I��U'$�m9)y.�(\ �9��3@3g�������#i�a��eU6_yU���v{z�� UZ�O��u# �Ȝ�з�i��i2���\�~XI��e^)�$<O�P�gu���ʌ����j?FԃUfY����L�5xO���$�v� �X֍:��h�3;��"�%o� ��c- ���ZhtM$�HX�d����i�kM�0�Q���ޑ�M/Y�w��R�~�x�}���ލ����~G�_���2<��i��4��*�����$���(�c���P�����}�0n��}��v'��`�P���A�L�~��C�V�	�KS��z�k���&�t����Oh���G�������PEi��?(+h��y�>$�W�~�i�N����n�Y���->8x�Ǎj��^���K�(�NxP���y��[�u&��S���馣|ByC�����/ �T�*���Z�E�0��W�۲�c�;�)��yN�B�Z,�v �1�O���i�O��"�����ͬ�	�?�<��cS����4�Ӧ�k%��l�n��k������lZ3W�d}�Ư`�F�tΎ���̆��9�zH�|i�Ka���$��G.����Ψ��V��\��޳��B�$R.��a�dߐ�"��ߤ� �OEÕ�#���.���f^JH-�p��G��lː���$J���s�������N�o�Ii�I7&���i�h�a{2��y<��K$r&���f�2v��#V��I5�|�����(IU3+�OV3"�1~A��Q�PS i$p����鉳���֯��|V� �������?�v�y+0X�PY��(�&V�ψ���Q֡V���˧�d_M�(�.�
Ҋ6��~�NG�ҝd�I���B��䗎.`��9��?����a� ���:��m���=��j�eq�B/��P����(5 ߣ����u]n\���n�i��̅��H�"m{��}`9�V�4c���*�]�K�H8U��D����
ͨ�,������?�7�5�.(��o���D�!9�.\�*�����'&K�i�*���(�Fe�Ia��]N13ݼ����~� ��]� fG��د]8��ϥj�ڸ� �C���WI(.jr�]���Ӑ�y