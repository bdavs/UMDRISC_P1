XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ӏ�6���"j�˿$��#��}�����`����4��P�D�80�i�����!�Fʧ�K�h֠w��:7l>�"S=_�����J&򕣧�Hte�g:�'�0����-����x����W�X�ī�)�P'WN�=��>S��9?v]��< B����^������t]���+k�6��ӷ�V0ڻC���i��8?��/�!�%��U�vZ`5R�=�;��xM&�m�F2/�l�	MDzw�X�VF�-�5"���žϫh����_��m6�;�Wֹ
e��V1����:����3AB����%4&�K#�ߌ�N6�?����[e�=�^2zP�Ù� ��-z릸p1)�	LOօ���.�$�>$.�#f#�� �0��F�JAbI,:`^eAV�̢g�I���5E�A��?[k?C���b�<Zڎx�����Lp�z���O/-�UX�q���� �w	��������,���.aV�+X��*>�͞�B��'���=B�&�r�@�����2�/�O�0[m;�&�Mʪn9k_M�����:hN�X%^���G���g��S��%*Ί
�����(a��EBP�&����nn�6��d�2c
������NY�w��˳�OzP��,����/
����<LK�OU�e��	u� �r$��	xT{�e���o��r�@�����^���|`�(�
&v��)A��G<��D�ICd��ɢ���;Tݟ���u�_�e4@�kyؤ�o�,j�&J��XlxVHYEB    fa00    19505����ɆՃ	���G�i�ܛ�+��g�*�){r���ч�-�W�P#ET��r��=�+��n]���y�|��]T��d��f�r��ADB�i�4|$�/S?�b��t�W�|��cF��=E� �;Q�Hx*�Ƒ��6ġ�-���#�BF��/�OgZe2Ȍ�dn�ƅ^�>|�+"��,"�y��k��G���X��fb�:Ccl� 
?g���Q��ɭ��ې��zp񉆷v'���d�Z/�UR��2���]�m�*�`lE���&Y�W�*���:ij�~�3�F���nӂJ!����c��o��,� ���C���ˌ�7X����s�u�����,k�W{�eƢ ���o�Zn��+�l�$��L4'v`%�ހB�
�N��(nK�Y)�-������Q]�f�O���h�E�B��k������;���W
X��J�g�H�Q~ػ4�ϓ�X�=��<�j.��b;y�^��C��SaJ�0-�_� ��B��/p	�U5��P�d���y�4���e�����6�nǆo�-(�Je��K:P��� $_Q�]D���q
5�
���V���5�;2�Ka���Ty��h��2,��c��c |lZ� ���4o�Ĝ}KC��z'&z�eK�;a�Ap�����$L ����_}&���7�Q@�zy����ߴ�g3�.Ńf�K�I��7-��r{r�zi�zv���/x�"�7l��|��4g=
� �P}	U0P����~I�f���/
��_1Q)���ʙ𳁹�K	�"���#��h���K����m��_R�[Z���d��#0w��_�UL�z	�qc��ao���+tn.{���8�h����i��2�x=tE~<9���|��V''Z`Ꮻo> 8p��b2�<��D�f��_x_Y3r�z��?/�m�zw�Ɓ+&֐��?��N����TŖe,/"Y,��f[F��������M���h4D��w:t��!_�m�Uc8c��F8v��f;nLH�a~1G���e��L��2sJ���i,�/���Zm#�u�p�fiT��+t�̭;��{�X�Z��Ie>�1g]&/8S�x���{_-�c�	D�t�����jox#�;�������s��}�tߏ�>�)��j>2Z��O��V��囿h� �Є��vu0���rC��[uj��^)�{q{��(�P;��a��RH
*����-����U�ӽ��42~�O&�h�}���"�ŏA-�Clv�#�1��T2�c���8H��A�t��U���|&wX��N�!�!�4�Bǩ�62��/8�Q��dR�]Y�Q�O��M<`8�5XG��6q�Y��W/RĒ9�Ēg�\tޢ��)'J/��u��1��˂e�Se��=M���7�|5��~!D�&1s�%��>l����U���f@i�����ՒR~�)Y_)s� j�������T�����6s�g3z>�"/t�%hd��m���b?\�X�r�����Y��٘8�i��{��I��v4f�)(�Q��f�u��&�� "V�h�{z$���$L����4 Q��J�<�m)��U�]�W�~�����y����A�?�����jpѠ�&oH����dG�,����ċ�7X�5GzΎ��px�y���q�G͵-,��5x�E�#@nrF�<)p�΂�DHl�,R��Q\���h@ P�3�o=��
-aF�되Vc2(?_�zl�NǠ�< ����tܡޞ>\p���'r�5���@�Z�_��L��t��]7�X�*�k}�TF��A:_Q��QX��r�32�f���_�l�Z���R��W��ᮈ~����(\�[��h'�E$l}�Ksy�v�?Qz뱸�z��o�Q��W&�\�� ��8&2os�ֻ �7�� �2�ܜ7�s�%�6n�ߘ$��E�:��v���pL�G;vf+/s�W�g����N��6DCie���*���s�6��i��'V��� w:kD�F��lq���o�_�jw�4!���3Y�w�@?!T}���v5��"�L��U>WŃ�\�x!⾒��ǟ��N�VOk%(ـ�+���W��s�Ü6���uj<�8�9S�4�L~����ʍ��HqǤsƥ����vf��/k������G:̢��8_�������hU��6ty��ء���"��n���S�s�*�)�+/"����vՁ|���ڎO6��	��m���؞�6,ZGNў/o�-��6:g�Oyr��t���t�[֚�Kjd�̷��h�oL,����w��sp�lr��>�C��ZN�d�	ŦZ�}��&4W�� ���Q�h9�eP7|"�y�1[8�JN�γ�A��4�	�G�u"A��p�H��x�m�L�Ŝ`
��E��Ff��W�*ݽ&�/i�4�LN+���es�i����b:����l�6��GA!B�g��a*�4�C�*GsE��h�N��Rϖ?�RqRSX�$���k��&<~#���ʮ�uh�K�A-�����k���A���6z�vk���6j6;�t]T`��$�a�@�Q֌)V�2��h���/��.�gDZ���SnvP;��
^�I{x�A��rM�)���f��3���72z�R�M>X V!p��[��M�[�A	[�*8�h�vY��F�"�7��9���A%�v�렛��s���^8��tCKv�~��fJ6�|��3Cv3����������^����@F�a��ݗ���b��M��|l�=��_���E{:��J`e�%2;�g�j֗0=F1�C|��L����@m�������pV�6�O��}A���Y&��y�����=�Sjs'�#������p�#`����0-��e�*F\�Џ��g��g2������]#�OK��:|Y���
��ǀ�w���0+��B3�?��]��c�Io��X�|�zՀ��Ye���uAؑ��F�K���Z�ɮU� ް�Pn��f*z�*����u|�%n�Zj/n��P�ro(� �y�9~t/�)��qCB�H�n���qq ��
�Eq9�&��^}��߯V�4u�⎎�b���x 9c�� N���4�В��QW�e�,07=��ے�2�Af9�-���S����MƸ�H��	UB9ɦ��i����^�o_���.�=\��a���˗j�	��Y��5)	[�L��ķ�ҚA�4����ߢY(��8�Hn�z�T��?�l����,��!/̻�r��Z�Z�:�c�{��jji�ns����Q���D���夽%yt(&���R��d���*��|���kVb�eш�/���C�?m�m���vՁ
�v^���Cw�d3�:z��&zoJ,x{�޻d:\�M ���9o�k��M@�[CK�����U�ǒڿ@����"���vu�x;��9k�[TU����#��	(n\ͧ��m�Z��A�����V���E�!�!�6�����{�$�>[��0ƕ;-�c�q����y���3���Ԟ�H���=�����->��v���4꒰�˫�~���eMf�ᆿ��Ɲ�e=EK���1�'Q�E�ѝѪ�s�*d+Q�oc��Wb�j����F��Y 9g�g�!��1�t�E�̅�ݓ��
#�T�r����r��z���Y#.�a�!Kv��,;3��uȮ�o���d s5da6d��4Z�e+m嘀An�|F�Uo�맂��Y���-�o���XyL)����6�����r�T����ݣy�� ]��!�.9��6�čí�+os�Z�ܯ�2үţ���� ^��o�[i���xb6�Q�iiKն��0v������ |QUw�
cu�dF;�R~vi���ԭ��4�u������&D/�F�x+�g�U1h�ܙP����q_m��ԣ�[H�&����r_��B
��� �zF§�XT������>���O&Z��E��%ϴF�a���v��
b?���CW��I�&T�q�mU;�D��/�����V*��O��}WI,�"�e��]����L�XGw+r�P�r�v�����т��8�� �ǐ(���yQ���*Y��P le4�W'��0���W[X6�����ȴ��+�٨�f�y������.0��B����aخ+�>/����˽��^hZ�M����{�0��� ]�LҎ�A<��`Ϧ3��1�Z�"D�9&�Y����X�'�}�cWh�R�h��#}WjTGN�s}����E��f��}�{�/?3����J��.5�������#�(ޚ��K*>g�B�Їd7�O�xP���1R� ��R��p`s�er?S����)�Ƥ������KT�O�_u�)R��w�����AH�A.i�*��� �&F��nn�cix���ZAIrG1�4�i�c'�����m�M�b�r��u`\k�ć���S�f��DTWC"�aU�*L�E����*���U2�b���f/x� �T T���$�H������i�ה����_�{�yԑ��dBwT��3L6�Z0�B��u����nmB*����=`��!���1��=�t���v����"������	��*�1�ѹ^��/	��B�B^U�i �,+��p�x������ğ�q���r�wMc�����jG���c����Cq�-�ø�bIA�����l�s�p���;�#X��g��Fp��q��4@+�X9Һ����.������M�'T
K/�ċ�v�����/�0��N�L��ñ��u)X=���� ���QyE�i�7ͤ8DB��y�Y#�|�aFl-�� ��eg������)����EH����K�?CS�! A.7,���ɐ,�?R0š��;���I�Z�z�$d�"9�1�D:R��v���Z>��]�����r�;O���\���ԧܘ�k��[c�/[R:'��RH�p��*��6CxS;�R�$Ԑ�7n�2!vja�����l*�&U�X�Y6E����<��5z)����~�^u�jA��C�zvA�;�*�~ҠH�쑬/�6%v�I۰���ٕ���~h�Sh���&إx��
��,�AK�*�
+xOK~�հ�G�4�g���{��0��8(�FVFds����n^���Տo"�X�+A!�6~m�*}O���4ڇV��±v�Ҋ��]��qJEC��i���`��ݱ%�Ӛ=���'���J�H�͏������B��o�+���^,w�gXw=�����.�R>[���u�jή)�l&���\�%!Q��H�җİ��� �=���5��0�wa�Zg��X�H5�5h2m/���`Ou۱����Ń=�gUe������h-�T*u��(���x�PY��&�?��e�>�ƃѷ���
��ĩ�5,�Bt-�~�M�H3�U(�V��)���6xV��9�n�Ӿ�=���3�	��ص���"����-�I���S"�#����S5���#[�Yٸ6y�5F��ɄgwЛ7���%k����Xb�r�鈙��E�xt����AM�WH�9}��i0[�w�^� ��]�Q]<�@�_���|��2+4���!<?�{�R��7�?.�����Ġ?P��hW|�0����A�����Ί��	%W���>�p�5	�'%F'�-��v�P��3�|��GE?7d���r���_Tm��x��N֜��L�B�,�����-B]����s'�s�.�B��"�K���trE\7�1#��kO�6NMF�O����z��c�-�&Ր_�Ÿ���W�T�c���n[#�S������[�1�\��AD��d�OU��-/'i�;���`��X�r�3'�d���̚��SӼ������":LL¨X��>�c7-�u��(��JQ���=
�J2.��bz��D��J��;Y��Lg4�Q^4z�5�}P l+i��Mƃ6�zJPX����aqk�Ͳ��R��<��D���~��8�J�&�mdZ�X��\.�ٚw�������_9��"Vܝ{�)\2�F��C��3�sk��6ɟ'��<z)X�XE^��p�����&�qP�o��V�ygҲM��[G�S&[�����%��r� 5��s7U b�Q�d�� c�1s��YW9}Zx\G��-4t��5
���+�E+@�4\����Kǭj�gc[}>7�Sʛ�]���q����5�XI��b����6�0���Y(�8RXD!�t���ӫ�'1M��;@e*35|�O�wr�mL8�#���sR��~iz eޔ$8��h���0��ڨް�}*�2�?�Hn��ӹS3��{G��d����e�Ae�`m`1�tYQTi���|8���3RS{劘XlxVHYEB    fa00     700ʜ[=���ʢ/
��:���x.z2/*�S`���"��+qz��d���Ц|`�sdECp���k;F��b6�+��j�+������B��-���%l��$��������+��-��|�Lk�7�^4��w��N�@$o׻�o��R�c�Y��ͷ��"�	C�fĔ��̴�YH�[������|�}��C�V2��:K��\	�IߑK�9q�t�����ʤ��^k\ �d������y��F���['��J_��H!e��uV(����\끣ߝ*���F�C#9cd�[����%�b���b�����L���[Kc�}I�Wa^�S0P�Oz�:	�5�7Ç|�1��8;q2;d���"��s�=Fi��i|��H��<��X�^Lo#D�q b����{��Cn��0�N����iN��#©�i٬K��~�r�6U����xX���@�B�9�u��_T�к�gՁ~ڒ
��ݼ"��n$a�\%����<��+��_�r�\�~�R�͵�;�1��N\#F���"�>��F+�G;v���MJ��\��	���%!��8e]=�8De籧��{��=Ea��@��ɋqb�T��͓�rx�ͷhR��
pyC�^i�û�Q.>;Ќ m%����j�M���3������%�����i_񚢬m�V�o�]���ـ�MI�Ҹνy��=:�r�!��*�̂X�mߤ:�|�E8_���T����F齡K���ۿ{	M�&���o��Z�3!s��j�t�
��� �˾�,�6�m�%p"əA�d�~A��pC1x��x
8�o!Bl>����(�	�;T?�ec�f�Z�%⇙�w+��Nie�g�~����bw�0D��[.:R���~���hrn���y��;(@�v�T��0�iJ��f#Y�c4�rra�T�ҥ
/;c�M�	�d���<�)S+��l�
��O�����d�4����66��2�غ�3��]
y��H�����_c�3��j-��0��+�>�zfXC����򀡺�iJ�j�@���X�=ɦ�����;�â�� L۴ˮ���D`�\�ܿ��u�fm�Y���ZuBpѓ�_�] H����I�3-~5ǁ&9��m�����~�'ƞd����1����3�F��Wj`y�+���d0r /)(�5�bK�\h�Q�?5����3��-��T��r�<��衚��&H]#ГDr��?<�E�W`ϳv4���>�kRM]�G7�Ťb�a�/.3]���^�_�ѱk�\~�"���G>�n0�@���*��Ɏk8�B�T��s��P=�o-f^N/1��e�J�����m%�.��M�YLEp���Z �u�����'��y*H�>	*�����[�Kc5�=:T"�:+�<5�!�1�d��/�Z�7��v��pa��X[u�����c���Ҍ�]�8;hɨ�U�}���H+�0f�O\�@�C�r����e��oma	��b*jN>��x�u�ݹ&�ڗY8J��7_�yH;��ri��:�5��5��;o0q����)�m �}�A�0�,��{�� ��}t�͋��e��!b�� �Y�9�r|���� ��w��(:5w�*n�}�^Ԅ��vR�t�$,��My���h<;��[{�ŹAM��I�T�OzG pu<����k�JǪb��M�V��x�} 0<��׼{W�Y���{���Y��:��/�	���/�O��[x��
��
bu�&l�.�fp.F%����e�XlxVHYEB    77da     a60=|	�0�ug�#qq֮�CII�X���%����~g?�'�m�����b�f��w,��F�˾
q<����Mp��-�_��i���]1?M8D�ԣ�8��$\㸺]ױ�k/�6x6}���zGd��mՖ
b�Q�T]�R�3(�+����m�ϙ۔�	�����8���?�f�tT,����(޲�V�B��7P��T�"�k.x���^D���)*�6Ր=�ö��:I=ζ��t�(�+ԏ>eG\@	���f~�l���E�����Ւ�wUps;%�sNѺ-�%��Ul�!�.F���>�EW��V��C�l��E�3����鳍L��m����{�;yH�dHY-�$�p"V�O�x��c�u	0C�K�������CQ���M4���S���Au&��>�R4\k����d���Vy�H<��u�/�Vh&�;x2'��z��<{����?p1X�|!djE��#��x~�P<�P��z�b��.��Ky�]I	e<C���wC�%愩�_�ܿ{��o)B�&>���g�~��ҧɊ�p� yi��@�;�T9�%RI5����2�����O84	���&j�Nw�!�b⤫�,�J]E_!�� m$��z���ϣ���Q	���ϔ� Bq�?�h����8�Z2��}j�����=���z�`V�S0�%��&��E���i�m�Ccl� O��V�.p1D���һ�C����@��9���o~�J+QAdd�e�ӑ���em�G��z}�������9��Pb`�}0��P�ZH��_��I���/��V�֓s�d���Սrx��u&��}��YMjc��C�
���9n�,/��̐V@��Ac��n���`��v�2ۂ�sb�E�"jP�~���a�?I�B�L>��Ǧe!>�+j]&+u��00El`]�R`�.�2�^͉�ph�)<|2�\��ayl�=~��~x38P��D:���'��܇��C���jT
�V�K�"�R
q�	EA%��^Τ
���ʄ�H��l�t�J[����gn�̌`rSӯi9p>5Wr�Y��g�uC�N;�����~[��NM�d�� ����X��`\&@ �BB\G�cp�O�=�ň���yE+�=�F�0E-uԃ�W�b����ȇ+�?�/�q�5��6(,o�bP��*:Yr�xjk5��,��*�ʾ��yc},�^v�8r����z{�UE�
s�iF�Y�[B֝���9���^��A9n��a�;ܐ}�s���Z�c(��"Bݎ����b��3��g�5�^>,�@qG���/�#t��zv�����m?Hʪ���� @£*�ξ!2���<�No}W��X��yC�^���용�e>o�?<伮ֻ"��V��)�ب���_��(���'g>��s�Ϛ������e�u����ة�NB�;�ѵ7\>��_-<Ɵ?6S���sv�
ք�(UP�U���A�M�?��z3fbUj�-

@��.�ݹ�[X�� S�%7�	�,�zB~f^�p�V@ꋢ�P��\�Rc�'woc|�/���}r$
�0�w�!4�^�1dh2G������A�1��p[QGe0Wq�H��Bp�eghMH�@��������w�:⒢Eϕ�ey'��uW]j&�r�3g\��3"���p��Bԏ�(`�^����h�$�'�����N+�[���~x^KM��(["ռ~�E>��d�0�!?�]	Wp�R(������Un=�4�=PJ1�q#1	�Ϛ�۠� qջV�{D�uմ@���S���%!�k4�>���k⦘�ff�%�Y�ܧې���s��/��(��%$̃�`ɉ�1��U!>-��Hd.�dW�=�}�	�2)��:��1��B�i�	%��燃�,��P����^�]�/$J����I�A�yP;���v�>aʮ��;��[#����j�����s\��i{�������!(��!h��e���F0I0�h$���M�n��KI��`p��Y�e�*iw!� �nF>Z�$���xa�8�1�9�*�Z�C��<�BO�IY��/��ӵ�G~+���O`�����qٳ�AP�t3F��m �A��׶������R��ѥ��\#��>�z�5�pH£J��	���*/��_5��=z���q!_ar��eg�Ѽ�o�:dk�%,��BDH�D=2���2�d����Ѝ 5Z�v��\�ތ��#���Vͩ^X�<X�H����_>K����;	($H`ZN���,7z��hU��}�G��Pg�TE�څ��~6P .�t\�̓8+�>�a5x���J.������]�� �?�i]�	�gL�Jx6�`M�J�R�B�Eᑐ��*���nD*�{O�?([(0��ǽ���9h��c{l=(�������`nm��k��3Ê獲ԇ0�������vԷ�(b�9nA^�i��O���5)�\2�Ĩ��
��Xy�ٰ�s����U+�&n2�����l�[�-5[��FĘ��耪�:���2����Wj�a�N^�k.	s���AII��"��	0��oܼBՅM�+��$ \��T��#8�ȁ��YM���s64)\Խ�ؼ�N�j̪��gd ��>I���:�"X�!V_>6&��7�