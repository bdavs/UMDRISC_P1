XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�G&4ِ�e��a(�2�x:ywvL�iT���<��3��;ɖr=m�b �T *�j��L�&�+7����y�?Ȁ���؋�����6xc�IZ[^�Jޯ�H��"mYU��"!���[��v�k8�΄�yN�6��F�w�)�A*2W��ۙ[,�� ?��Ȣ����"�vJ��:e�N�3�S��lG=�{#Z�T�w��˜��yΘ����U�z(�3 M��%�<�NS�0��No��W�9j J�7��,ϴ穑f -������X�Si2�i"�����2��%6�;]^�W����W�sWo�l\A�R����FE��V0�F-�j�y*��m�t<;���;ִ%��`��*�;�*�"R���c��e�	���f<	����".�~�Ƹ2���9�TǙi�-���t|�q������g�����"C�O4y���[����x{�W����@�/uw�<�������
mW:�(���
���qb�JdCuh�����(9��n֫�=�	�P�O���$�@0+ �	룲n������q?F�A����4�?� Ml%�#Jg#�)A!��xsc��g�9�lkeA��,���,��8@�҆�R�D__>ig!���/W�콋G��,&�H9�W��a�,L����S�PU�A8������8�x�p���Љ����xIa�S��
9CD%{m��[�`�~؛�B|�`^Vu7q���d�f��*�8%`�����U�֤:�����LVߋ(��4YXlxVHYEB    33bd     c90 �0/�<�o7/�����W��w�q���"Yw��]��]�.&��,%�L�v��"䯲1��S�����Ywy=�`q��<�P���J,5���NF�q���;�&O�,�����1�L������5y���v�����4��&�#�Ҷ����죔��F�I:�2!�����o�ֶ̈́ _������y�бg�F��-�v���}޷�sIQ>�K]�0��P>�Q)<�E ��������Z�.���]�L�\�S�k��&���A@���S�����;LШ"����i�qɗ�$|��DM�Q#j?4F�XzT�p����w�@�.� ���f�@'�p��K_��7��ts�1��q)�����Z�t�����~}s�@�l S��?��S�{]��Iw���Q�5U�#��� _ç�<3S�t_3ϫ���D���+k|	:Ơ���K���I�׬[`y��&S@�m�u��	1�BH��YVD�X�Ǒk��8~РnɽP�Bu�Η7_���h�6L}A�qEb	�6x+)o�M�n&�ql��$�g��`��[Ȩ.�/rt��vb��avjl�ˆ2S��)�V=�|)��V�i�5ԙm	�<�K�^ma����x˴�P��ΚqM~�T33�(��{�Txj$r��?�ո5�E��w$�wO�;NGb�q?.���������:��=��$��R��_�c8]��8��Yh�䖺�#�Ol؊B��/�xg�3�#L��j������)+~H����pe��]~�;�a�zvG������]%5OV�7uT;W�<�����@cD6�ƑxT�@�,�6|�C�
H��?r�\wU�6�4�6����Ă44�G0q�"���r��b�J�6s�p$�8�j��,�.I=�	�Uv3G��������]3�3���t�)�KW���ԃsv[@�F�v���85��������,F���Qw��h&fÀ�6x�,�"~'0��"��U4�ӂ�]�̃�� �ڍ���������o�xS�:]P�z�����깼�u˘f͌�9E�;�7#�+9[஫]�����P�+��AD(���6�r��r��ft��o�F`���L���~8�ܓ��BRZ����e5+Z�b�[?�+���~��./7K��B�^��}I����/l7���׫,���I
7[���cfe؄�e��<�R꭮ⳟu\�rgd�4����\�p`f�ı���P�$)lm���7?�?�W��A�'S��>
�Wcz��Q��Q[�<
9���~�8	��MY', E�坛�1�r7�MN�(r�0e�3�Mn��w�s�$ڰ</��5Ie*4}�-��q�p�
����j
�ȶ���,�<,9}
-B�m�e��\0�-/�p�ōc���|�� �M�t��Yv��kU�����}:G�*��#s��[U���t1�G��Y� ��.l��bW��L(7�U��r�q��c�'G7%uY�������Y�|B63��k��\��������Ǝ�VV��NX��r��#�Ә�t�)ܗ�o"��t#s�H'���q��������R���WEel��nPp+�t�I����LB�Ū3��9b5Gmp��W��/�����j�>�q��������К��2U���R�r{dsw8��4
�Mȕ+A&���ܫ��f��;�O~AQ�������ٰ����q,.h.����7�ek'o��l��,V���S��4��B��$��|���D�N�Ȝd����d�=���>�g����ۯ9?�hE��Y�`C���7��)f��*v�N2k��O�@����Ksc�#<I�%tW�C�\����*A�%S�a�4�q�/5�ʎK&�2����F���dJ۬S�.�g���'͟�����w�J������s�i����{�\y��YS����Na\�fG�g�����R�Np�?W#cx�⯢�kO�||
�Vᓀ�>�Sz���{�ݳ�õ8�4�4�Ͽ�9J�I Ψ=�OK��Sr����9���;,�]�
��g!#7X޻�#�Y��h<���8>���[�+d�Kf{�:����^�e�2s��W��L2(�3Z����c�Q����?�EGN9a�o`:еŹX����r��M��A�ڲ򃽁�˄�X�§�7'��}|"����ټ��5�O��|��Z��S
���)j�F\�R|G�I�ӻ�;}cI}2�C������\��պ�ވ^Q~��Ziw�]�I�{����ϣ��*�����IXs�`Uu����a�Fxc�ip�0��,xa:�L��U�۱$�H%�io�A�@�a� ��M�_�LεD�%9�gb�=�����D��y�]���&�Ŕ��5���9:g.��>+�|OG1嚻G6j�@7�p��H�WY���QS4E�f��Ex�m���� �Is'�*���/P�(�}<���_�s?G��X� ���7B�n'�_��^����l>x�7��Vm(X��	)��?OL����l_�/&���T�`8��%�,�RmH�|s{C7k�P���ٗ�}UVld��Q �*��vv7��I��v-F�G�u��,��X�ZZ��:��0����լ_�|�9������D��{Ak�@Cy@�)n�즟ƃ4�C؍(�.}5�K���Sp@M|�R�n�X�פ�C����c�~̖*%xk�p�T��P�����𮲵DC��(�K��[�Ń$��$i�O�(ϱx2,�î��d"�>y��w6�?�aI�^��Y��N�?��Yؔ���Zԟ[R��Z��l�ceݹ=&P�"�����Zqʌ�E+�A+k@�Ʃ��%o50b���|�H�,t�n���]?�m6���P4[l;:z�*E~"#CK-~Á��R�[TF{��) =["��c�-�����&~ĝ�#E9�ȳ%��j�t�<�6J�8r���G`QL҈���04/��@wlY���	0;P����&�t��Z��qc��]ᓐV���·�J�6Y.m��sB� �hX�<��tH(@>A��IKS�֮��O�2�[����w�,�uV<���X��A��#�������L��I��.m�4=?LvQ:���Ff!��0��"����1a\�����O�N���1Xq�/��&��"�Ϣ��'��s��n���mb���p�`�BD��sER%