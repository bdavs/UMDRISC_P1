XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Rﰲ�
p&%7c���I�)j
��E��(������
χ�.&� �L��[�7�J�ҧ�u�2���G����p�?��J�hW@n������)�����m�9�_M�G&����Jf���~3���rКs�1��CT�����-�= j�� ǽ�����t�(q�s��R=3/0�g&q͓ �X��:5�=�,ɘ�Ή����t��� �K��0��mQ��a�(
_�-?�0і�겮k*,�<�6u;F��_�l��}Q;������H+��U�9i���[\y�lC�D�r��o�,�@_���e��묚!��ߞ�)2n�R�Wn$��G���36(���T��}1�����Vd�i�N�̂F����_��@�i_E����y��?a�S,ûs����=Nb��&����U
>�y�6�����Ҵ�VO��Z�B�Nz�c���X�,��-]�$�:|e
Qf�E�@Z���v-6ry%���|��^��2�3I���Y���
\ug�K��6��[�ʮ|�w���6w7+ʺ���y�J @���@��A�~T�n��|�Z�/��䜺T��#O� �r�%�`n�8qTQ�qã@�폜��,�$��w�*y�a,p&z%16yw�1f�������r�Y���r��t�d�틵�j ����¨Q��~�r�����4?i�w�D_ӼV�9%L5��Ӓ2d+X?�ZS� ~�'���J�z��==�Z��?t���.dbB��8��i�Q�:DQ��XlxVHYEB    9de1    1670�X.S�����-�-#��F�9k��P͓n�Aɏ9���}��%�GP��r�7����0�����砺e�\����%Y���[�L& �!�G��!IrY.� �#��Ѡ������S�	�������(�`<�ޭ7���J(�|�{ �(b��B�C��`ѵ���(}�g������j/`z�,^���}u6�m�li�+�"�eH؃���N}��'��B�����Y�Y�)�I��3v�� ]p�������ߞR �Ԫ���w(�K\���tl�>t(mP���l�!.}�Mq����!�꘭l��տ�	��,6�?1d �p?(��,FcC~/������ߎ�_�j�a���lF�q�7E1�y����@�Q]A�=��#��_��g�eEɲ��w2/i�E���|�^�����_ q���}E�!`uR~	nasUv�\Z��0�|��\%Lk�7�,�����U��њx�>_���tj�����^�Z}��'v�אH8<T�R�1����=������w�|B��"�k��G�Y1�Y���(u2}@?�o�l����S������Rl,�I���,�1֋�>,s�HuxR�]u�L*�=ն�>e�J�ߖY������/z ���P;�Y��ǎ�U�IN˛"��䌊��}d�C�ݙlX.6=Ч�f��ъh�X�q,6�[��ϩ�U&�;���`7�z Y���ь����ƌ�~gN��e��È6�mʎW�a��%��0�"�Vi<o#uh���5�y�`�k����X�H/��1�M=���P��~��(�d��A��r�ԥ:���<6*�Ԣ1�A"�z���5{��6��S0�*1�H6���}�C�!�ڀ �V�۬����K79�T�kMGf���mK�g�ݓzwE$We���n���;Sή�{�+�4d�#q����	�E�<�+.�U; ��A���r*���v)]0wl0��Qo�>?h3:�} ��������%��T*eo`%3D�/!����4#n7p�-�PN<��*PN���@�/k/k��_M|s_8�	e�Hf��^��ۗ��F6j�R.��g�o�@�ͅ+���8�a_!��D�����%�V�y��D7���`��$����.zy.��^�n��>����H@�9����*�����3��� ���%Lz�5x�m��Em�/�G�o���;��v�Rp��h�t�s��ifu(���/֗H�a���M�:�("��t�viUל����?�N���"2�x�`�������,��g|u�bb�MT�[��<Ah��0ҙ|H���F2uZ�4��cbz����� �%#% 0�&��OsVڌ�DXdU��� i��q���o�"{����W����)17�y���~[]��I{"F�L\,�������IṾ3f�/o����Rr�d�i�9�ʪ2Z8{�	������6ha +?u����^�FD�:��UTu�����yS����}���4�Q4�_ߔ�'��(vY"����,�a��3B��*4��"z��{�D7�uK�wiPIs­ �ů��:����*�y�k��/���\΁����މ����\�;���_��H�@>="�8�L@	䅿=��C���]�}S�i�i��vY��[���B;���B� tҋo0��:`�z��$z��=��WS*
����c�
>k5�-�Bt-�(a�d}L��d"�lߨ��]���������#f�[J����B�k��ʔ�s�'�/z�F��7c*ea�u ���#��v�u4-
,u	��m�A�ރH�?Y��g2�B�&�+��?��I~�*�\v����ib~���٫��$�\��!l�f�[�.��|h1�F�D}"6�.���r_0[Ջ#�:�O�(�W&v�f"z�X5#5V��*�W���G}�A�+�;�#�]wz6�z�FA{�� �M����
w�v�:���1u�'	6���ew�ɪ�5�j��{�g������t�Y�ܕ�����������t���q��@�I����7j�˳
��͑q>a
E.�h��SOr	>Ř������Dp�إ\�����,��2�I������jNԓ {q��yi��>�k�b?��!L�=����He�_?e����w}�n��o��X�=;�XQ8υ?��v��(z{bY�d���(ȽGx�d !�D��Z�p�<��:Hg�.ֱ�^GS�����_�����0�v���3+hw�D,���C�XL�����Z$#�,4�lT�Փ?���Ef��7���|r'�����85MLv%���}�!M	�TG�U���b:Qxj4��.���57\�%��69ښR�mˑ��a�^��i�<i`�te�����nail���ȏ�) �v��tBa6w�V7�YV��|��6��&i�{�$�:�
�Y[B��WL�����XD=�f��2�]�u?5���^���$���kז|;5*f�e���Hz�����T�MF0�)�d�Lt���� PPJ�\L�S.�
���i��m�*��'ol��Q0k+7/�Y�r^G���$��pN�ڈ��\�x�> ���T�@�!ׯ|�԰�Sk��"vv{�*O�0:@\�NrݺYc=�bO�Ͼ�Q48k���ϊ5�c\&L	������w1 � �z)<@t��8s-��G�I�%5^�4�f�Pc��1�L�kq-��F�
WQ��	�܅%�	��TCZcE'�H	G�f*��gcQ��R����h����
��jw)�+O��}E�!��4���	���Q��O#�S`!�By!��͞�\�X:���e���'q��̴1�xF0� �'>66���)����N}��Tw[ew�-諦Jaکzﬧ���Wz��o�R�3�|%8�t�+:�D���/��i:���O�o{+�F�g��6�sگ�X+��g�{oO����?��:C���*�!���e�g�)i+)#����t<X��N��Mb�����'m����
[�qE�K�]�cp�0B�2]�x;�v�,�h�nۯ��e������fE^ºȅFۥ�����60���!��d��ٱ̔/E��(w�W(b�	�Ggtؙb��;��b��3�֗�k����znR3,�A��N����J��������7С^�ʃX����T���30Og� � ����1*şҒ�Qp}"6L3p�Ȯ��s��\�/0W�^�{,�_���QX��ٽ:�h���W&�XH}N��;.  q*���
�X�Se_�|HٙH�3��<�o��������:�k�h�sy��g�ǲ6��u�w3^c3�K+D:j��|r3,1�V���{�QYw�20�D�+�X���t"8��q2�)ׁ�.���FԞ�#Z��P�>�3n
�0���˶�{2�7:$�$��&�/��p}��\<$�<̨�#���Ͷ1��C�~3o��҇~@<]�������v��\H�xN�w�xi�C$�R��u��m�,-l������dW���e��TB���TЭ3�L��N֚wuH�t���ؐ�ǵ	��f+Q�i�X���>�V����|n���+����O��1\:�z��1��33@~���ILg;N
���s�{S�jr7�C�TP��O�ʬ�L�����(z0泗�C�G�Tjc�bϛL���3��_��l�v���u� ��o��|�ñm� K.���#����!����2����w`�ﭱݸ���~i�0��w�?�����U6Qo�p�W)��>��5xnUD��f�>�@��'�"��k�l��h����uĲ�⺼�BJ����ۅ�S V'��e܏z��	��I�p�����an@rqa�Бp,���i�0��%<f����F�{´^����ߕ�rMu]w<SV��&wBB��U���{m1�u(��ME`�z��.cSi���?9��h\K�M"#W���0�s0qeḪJ�˞e��iƏ�EM�LV�����111�g�H��C�yv���[��< �/��� �oZS��Vq�����wܝ�.;p��@#��7A �F��`�|�yny�^�6/�i%�L[��/'��a\�������[�𹥞>���x�֏;��&�o���΍M����e{��Q��S2��&��[�a�����W;[�N�7�-Ɲ!�nF5���� )��nS=bS�9�z"�'&
9�����uF�֑�L☊�^8[Se����e��l"COwѨ.i>�`�I5�(xz`;439�u�=��G��8���,����q�P�ے4s%�E������G��� �ЩW�oH6��Y����3$�`�y�i�d�|u �K�T@�͠�.ZH��!���������Ѽn3��`5��]E6�%���c̈́��.c�:�����ҁ'Ps�~����k�M6*����*�0����]&�?+��?Ͽ1�a������g�G�*xw:���
�X���V��k�]ԱER.�j����V�2�ǒ��ڸ��6��^'���u��.C ���H5o���p�]�V%���宕���	����b����fSU�~=���&��V�Y1��u#K8-'�B��'w�6�S��${��R"|V�Ё�,��=L�A�_���̂۶�}dQ�=�O�k�qt=�0ʠ�1�ƿ߯������<��.T���!��H���K���u	��G5����L-���20b��/��V&�|��/X�6Șr��:�MC���w����ʟ�'��3i�j�'�2R����I��T$�2��:N��j;�����-C��>�����[=����pV�$,	�� ������O�]�}������ι�uƙp <�?�`g���6c iXm�%9���"��s@�Z����p�bZ�����j�L�������&��GD�#W�*a�2:��v�~7��P�Lɷr��%��֢��G.��frTVf"E�쐠~%��iѰS�m�qġ#J�U~�Zcm *;4�n�����c̽ŘI3�=���g��5W�c�m���;��S�C�����B{B ��w^�3��[*�Il���F��&F��W&?��ෟ�09����������3���)���u(T����}�����A3�Rt��ui�z���/!�B��Q�~yh�o���ԇWZլ���j��-��:%ԗ����L$��=���S5���ҥ��Q@�ĺWi���6�y�[��0�'��sȉo$���@>k��|s$':gOVߕ�Ko� ��c`}��J4uD��9��Ʃr/IͲ��o�%YznDޠo�>&��
���#������y�Ӌ�@MG�S4oqE4���wV�>�"G�����zm��@��y\�Ʃ�Z�۶�*Lqq��lT�Jd�ɓ�N !���QC���0��(1M�j�d{��ǂ�G����%$�u�d��U��4E�u�
�?u���\5�ls�"� �2���6��O�v,�� ��iY �	W�6%���”�A�[�Nǖ�$�by��ƌ�C�,�K�Be�_���� ��|:�^|@Ϸ�c�k(�Z��XQ�C����Y�Y���m4ZX3�k-P����V���0�\ Qmc��j6,��r?�\��F�մ��9<G������a�F�&����L>`�:�PD�؆���b!'�V�Y�������