XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��FUdh6;�9D���"���2��nl��%[K�[��|�>
�>����l����]�ҺR�~ܔ��hj��.��?E[@�UƿT�CG�y_d(4͟ ROٺb}�S˾�'j����������@!�����ێ`O�1�Rޖ-F�`�u?�1�۰  �9�+ϊo�d�#�[�UA%wV]�ʓ��2%���h>�m��T��>LcV+��ڔ!Ve{__�3���Y9uI��e���d�M��V�`�2�-Ƈ@<d�G̟ŮmU{v�O�e�X�ge^����:�.����-��1Z���W��;��m��0a�6:N��̹�k����� x��iV��1��<�(z��a��.WQ6��r�>!��X%�2�\�n�[f������T(�9+�����萖����%�. oz�eaZɪ�~�s����4`�õ}.�IR������Y�9fϾ���{q�*:k�W뽲P��T��(��7�j������Tq�.r�
�����!�F��|���e�z�D�tc�> ��M��O
���aï�1���I��FG;��in��REထ�`Đ��?�L��b�@�����^?+O(��G�,�l��E���GAW�]{���C��~�����6�6�W)���O�@�%b.q,�^�G!q���"@��4	�m|ʧ�^:���V�=��;�P�bN5�S�c%��Q�I�~�8�[����"����OxH3(K��}Y�Ǐ��-X���huM�2�BXlxVHYEB    aa31    1e409�ļ5'wY,z$R�%��H�ݔ�T��#q��=�=�{�]9����K1�*����!��N9����9`��g�Q8�c�b�7t���U�+�*�E�s7���@���d׭�sw�i�n:��
JK��ex,��YyV]�d�!���_$���;ؚ�кkE�C���y��(�J���iNꔭ	������0u�iї3vRx�6iki@��Q��d�7�ocZZr�봹���[
7$;����/~� t�k&�Q�Kq����D,?}���VqG����ßA ��<�ը��VA����|U<�2(�ɤ̈e4�FQ-V�L;��+m���Uy�K��՗q�Z88�?��u���� n�Lt/w�F� m����<M�=�������Tm�֮���� MԛU0����¹�|�C\��+ꗧ��5�#ap�T���NP�\�NDB��L�N2B6v��6��=�}��eE��+���J��m�j��*b���YK���`0���2�w��d�PGZ���M����Bu���n�����]q����d�z-)���	9�c�⛕�޺e?���iE���?����%-��Hs�YL��t�����Օ�L%
��������g�琢s}Z��� l�e�Z�(�y|��ӕ�8��SU^��h׋�m�U��ٮ��(�Y-��2G]��<x]�e��w�<����+`� ffΘm1I��t�(��z� ���m�\6
z�k�â6r$�
��z(���J����o����~������q�龗���<«��#�(U�#�QYc��4�$QQO�z4��3	�
��^��!Xru@3��zrS��n�3��R꛴�@��{.۲�oF�+@5�E�	a����"4����~��������@���t�b9x�UX6�:=�	�XdXRSt��A������|��w���<#�>�V��WDi�L��*��܏����{�F%ЕV �)n�h�3[Vƻ�X�aok\�����@���*4k�,��6J���$�	�Pd�\��!�Ju{�K�m�5��j�<�r�n����?C3�=��Y|�͹wlJ^I���HKd漓��{���D,Jm:'k�=o��`��m
�eS����T�f����3=�X�mi{�ێs��x�GS�u4H�v%	E�1z�T�4�#{����"��/s��1���WrW����ݰ"��{�\���C6���=�_��2� %��
��*��I�-S-�┬Ȇ;B��8+�NnQ�+
�wgF�c!�7�/'��(X�(����,��J�������K���_��*����7��qY�>�np<f	���<�����R��V+w�Ϟy��n� ț�;�����àX���'�vkl��=��-H��gK�hO)��|*Κ���ǳ�����,��*����I�+�x@�U���ʢ4B�$��V�_c��)���9=z>���zh6?��2��N\�hq�6x�c^����F.����7�W/�S��O�=��b�F��O���~a�i3>7v�t�����D��i~yR�2.�G㿅K����J�-��� �f�q�Ⱦ~B����K����S���Q����}C�7�a 
�����us����.ޙ�ьz����u-���f��/���r�wQ�G/�)\�+$�,}�1E"g2���@U�*�ȦDm :P`��m7�S��H+�\�%����k?s�Aa��E�n�]6�Li��M�I&���]etFXikDҏ��[��^at��n�P�О��B�X������Tλ��N�8[�;H?���+�f��2oBB����Ϭ��6�v�YA�ؘ�l��S�NS�*-Iy^h@0}/���KiF�T#�����!�J/���߬�����N�s/��N9p��6/��η���n�.�b�_?e�.��	Rc�N�+��t�q� ��X�5�c�h|qNžb`"f D�5\ل|%���^]��[��~vR{?��݋�6����I~��9���m����;R�*�d� ���<�XFc)^�ʴXh#���k1�JVi�<�{𹑨�IqJLgy2�Q��g
6 ��v[�ͲʩƬ6�8��l�s�Q��B����y���W��Ĕ����&Z�\ĵE�e���!�@�w	��d�h��j��|��F#,�sef��d���I�G66!C6�>vB�O���=�s/�A�_1�P�ôʹ~zW3|QF��F��,��J�o�R;�3���}�"�ŶxD���{~�!^;|����k9���%��~5�.�0�%�v��^�Ȃ�����U������ �?jľ�U�cG�K0�I����x_Č3_������֖�i���T�:���(����.�lO=�J2w��0?��I@�vz��+X��/3�~*]TF�d�������!�]f�u}8]�ǣ����r�r/%g`�������B󙹚]�W�~�c���N���:s�-+�IY��+=%]�/~�)3���s����p �(b X�����,���A���y��r�5g�c�=�>[�i���?d*����*�gP��<�oݶ�Ff�{j�T�X���������>6	�
��vC���M�_�'�36���C(C�x�N�s��E��1���$aw�HL��;�g�m�t�UU� �p���7��7=y-7�\an<r��_�/P����G�5l�o��H<I��qa�O�qf�M��?���oU�u�*��
r���\�C����}B��`��nxoES����{������ԧ��|��;y��j���m��rj�5����SJ�+�����a�=���K��:���q�ߡB���}���AH,a�"��vN�8��R�ڻ�YP6}Q�)d~ � �:�Ihy���b����љ���#��6��X`Lte: ᬬ^�z̊�O�Wu5�LW��ݱr����}9���T�6�$����u�?u��u)����$�G�K��*U��T�J+��g�`�����0N*d ȳi�(�C��h��芦ނ^@	��{{��<�O%�IIc��Q��y�Ua��!y��1�)�"H!"$x9!&1��?\ta�w�$�&�Y@"ڪߔ��6��uጜ%��E����M��f^fYq��h���7Hp<s���2H�S�ن	�p�<������L�O�(#�.���B)�ÇVmn���l�O��. Sz ���ْۗ-��#�A�w�.Y~� _�����U���	͂���u�]����݊?ev�m�KT�(��!&����p�g�-M���o,Zq�28���I Ɇ*��X���~�TF��4Rb�!�O��ni?�k#+v�ڜӝf �ڒF�~;�?W-w�<������:��>��w�x�[v�倅�S�f#�:1N�����U|�笸�k�h'_����C��������0��Os&�6�J���6�`��I3�!|[�w�	>棺��hMXoT%��W]����v�ɟ4�Q�W��L�ҥw*������6^C�=!��w+ju�H;���{�����=d)T����$X8�{u�v��kC	�%ߙm����U��o@���wۿ��� o|yE�ǫ�|�y��������y����~���۳IF��>�ޠ��Z�~��L�vb1E���ڻ;A�r�7(V-kU�%��x��o���z^4�+��/94�)�"\�ʑ�/�Pޔ�|:�����a�7�K���:����oM1�&���?���-lJ�5L&k�[|(�R��w���RǘtBJD'�=��vÇ��)�Z,:7	4<\Hĩ%n<�1�E�1��p�KpY4{=B=��N�����G�-�)Z�>e��IH�i���ꮽ���̑,�x1� G�y�j=��lv�!{�b��d�y6�֧*�^�?��Ȝ�ƑH{5�_�i4�`Ca��0����]��lA���vȭ�
h�7��^6�H](.h����,�ܴ��ނ�T�g���گ�-��T����i��X�e��vLd�d�;p X�:E�`�WL<-}z�.\������U��֒ p��ߗ�����^����=r�:!n]c�����7d�Kܠb1P�fu��җ��Tv�e��r��Ԑ�n;�M9E�B�H����1��@s���un�3�8�_�'������Ba>���2�Y9��|2�_�`^�&&�j=h��?'����1u¼���'��FJ�+UP�Ѭ��8�-��C��Ζ=�<�B�pݲ�qRi�^��hY�1f�J�Qw#H���5zF&��7����2f��K3�4��)��*vn��}V��r;��$<�L�� ��:j�v2���R�q!�,\�>�` �%�J�v��D���m�boؠ��Ig�����p=�@1PP��H匷�^+��&Tz�X�K�G������f��""�>��Cq��8��-9�]*<7F��s?���V�&q5���cZ{&]�y-.�A��0xw��``�@<EpY��	�BBՉD����9]�;���Y��%������!����h�l��KK��Ҹk[��y��Q�~�B��Y�E<�oO���`���pg�N�;Q(ACN�b�k����n>.�}xr@7�`h��y���.���	��<�xC*�����<�-�({�,������JC��\���y��;n��a���U]�@�X�T('b&��N&�ݞ�\�L(��t����x���A�K
9^~��P��[�Ѿ_�X����[έ1fg?/�C�hk�����Xյ��K,Q҄�����d��Z'����ۼ7Br�Zܜ(�x������ Tܜ�r��	�R`��z^���#r����V@�2��,�����'�Ey���>`�)[�Q,��u|'K��$\�Ϲ�w� ˄3�o�S̳���sR����TZ`*�A�d⟧�W!�S4�h��<Q���>[�{X\��P/P��YB�5T��<�x�,;��bq3o�+c���1�&�����]�rdɷ16K$��E�m~8�u*�7]�*���?�0N�&���?�SQ04��zUAҁ̠Q����F���cF:Da�Q�.W� 輮ɹ����y;��}�<&;��U2G�M��=��F��F��֞I���2`&A�,}�P�m5�;����ڏ�B)�YU��i����N[~˹�X`��w1��e�}�Xr�	w�PK���P�b+yfz�F�2����܈<��Դ����0��dA%|���e�i6�G���#Etb ��/��Q�_XR���rJ6�<=$�o�bi(�Pت�9�A���ek-�w15o�|̀	
��gpƀ2����U�-b��u�z��4]�m�>)�q���}�x:��g1=�7��@�S�J-��%�B:_r�p�ٯGiB���dw��26e9P=�1�`E���疺�O���Qu����Qs!q`4��Z�[< !!�&�p�c�\`�;XBOUs�f���R(C�m��W�e��y��}pI��^�m~Ӳ�'��ċ�)����?w[�ҝL0��p��y`��[���G�O�U�V�oЕ7�q��ˇ����\�r��]��X5J>1��s9������{���"߻��a��x{��&�l�� 6��Y�Yi�T������`|�p�漄����i��\d����/^�s�v��M���� �bMд##(��Q�5��f;��WA�1��X��5�ю���2� ^�#����4�ƶ��|N@����bG�W:9��i�91���:����=�Y3�@�{�ױh�Q�����[�X�皸#z��*\��^�&H�/����E�7K��w�90F��7���`˜�$;^c]��%6���E��O�+5�"&9������D}T"�]������h���o4P���U��N�W�G�JBYV�3'R�׼�"k�y����[����P&�K���!��%�9�ޤ�-P����Ӗ�b�9��;�AQXnR,��a�1�����xǃ�;�j\R�n-1"
 �d.^�D�)>׈O,�D���d��� P&�����KC�O��KXi_�SA��a0����0��|��v^�'l�D!vHsR��e3���0)����'�:��_vŦ9PLU� ���|��!��m��R,�V��gn�,�oa�S7)�7gp���T}�mL�ja8?��Q �zZ�	�����ο�E���t��TȮ���/��ʇG����������"�Aη7��2�<�	��Ɍ�.�5 Z7���s!��4�����%^K�a�@Ɏ���5N����:��rR$���8"��Nv��z�����>h9�ӻ*�8u:Y- ������{z�ϝ\v�D���	�/�)`q��<�!�(P���d�,m��c�i�=��	�\$M�֫@��'�Ot���ͅ��o�'l����L���ܳ�H�(�${��P��jV�h�]�6��{+�źd���a���Y����^�����z�E��K�� R��3���Y\��7�j�?���'u�e���?P]p���kA�T����0�'�������	�jڮ���:� ��3�'s�sH��E��I��IC��r]�Q�Z��T@I��Wcؖ�W��EM��C,��L
a����b�6X�$UB~R��S�� �p�����:����*YR_܊����QQ�[F?7����E�1�obe��/��x���լҜ�443��d��$J�$g뽁s�+���+żM�	�z�(<0 |}H\ј5��'wD-y���_�T�O�`�»wȟ�����_��A*iצ=�U�X����kY����X�t-i��vh�#z���M|h��u6o[�?6 �v�K�������r)S;��Y���?�����W�4NG�@:���rE=��JҤ�=T{5�w�I�����{�J۹l�����B!<]����E�+����D����̓�@*[%��ܮ`���^Tao��#XGs�a��3m�Pyya�B�����ѯL��_������}ƿ��N�5w+E!K�h��-�ө䞣�ZM��=nI��f��:.y=�6`ώ�ZY)���t�L�B]36���gWhD�F-���]��F.�o���Onv����� �M�de�ͣح/��gde���D�����[q�]���v��wS�H��u�����l$k������-�!~+�Ұ�ܸ��3����-P��>��v����ɞ�S �b��/-EE~�~?>JV�GC�}��J�ň���Z\���Վ�/C���E\:k���؜w��pgh������6uoW_�=1HK�o��I{���q�����Q�5&杻�b��t��A(���A���h��x`y��窠lA24�%�<<e��L�Y�����k'�5͋��WAu�I���]�s�s�"�<��C�z�:�Uj�.>R�4�m2)S1e�C�D&XA9�
1�%�_�Ci����p�saF!Ӌ�d��oy w��ͅ��V�f�ˬY��a�znQrC�|�K�)��Y�(��t��غ���ʹ�C	=ۏw�!j�d���B��=y� ����ԥg0�q�K�TF�mV��[��e�
G,/�I���do���*mKbL��P�hx���#��z���tJ�ږJ܂����HI8�݇�
�m��z�v7�m��