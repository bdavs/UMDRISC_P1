XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ⱥ"k��A�!��#��֏��E�{�]J<�����R6mD�*�%3�e�����>��[�hBcH.V| ���b�׏h��9��o���]�P�ͅ#�R?�<=�L9Jf.�TjD(�I�H�9�Ȇ�^�r �R� 
����@h�a8�W��`��?�W߽�P1p��G�Bs Zo�̶o�B۠*k}<]Ʉ���ʹ�G�x��м�����4GQ2-�/������'��`�9(f�&$I�W������)={�u�Bӈ�����@��@�,ҟ�Q��a0 #~$>֞u�j��I!�`:�7�;T�D������=)Ŗ0=��X6��k~luP�K��A��Y) �i,�q̔Q��6���J!C6��A?�5�s�h�A������fs���c	��7(�@C�Y�ı��m~C�43,�{��$�⼊+x�{S�y@���&|�ݮ�����*��f�*S,jҨ�I044�#�n��vծ��) �sߌr�B��B����ri%�\���~�+p༈iAB�]蕡w�w�iב�Kc"i�+�uX/o��~�Er�kU�݃2�܋���}UȐ��cg���DyvtG4C���.�����/-atD��4gϾ�eb�[�u�P�(09E�>�ק�Jc�^�u�ȉ�����+�a ���{/�/���Eb�qmo;�[�4�Y�T��h,�P�-��xC��4=1T��m�����r{qI�-6���t�i�F�#%�ChC����IG1XlxVHYEB    fa00    1fd0[Nc��t�eH�ְ�7��?e�o�`�Ƥ�S�����V���
����±�)9�Y��e��HA�M�]���zJ{^Yܓ&�
r�4�'���@TX �Y���,�\b�V$7HWb�6�G�h*��&��kW�"�ڱ�Ũg1���*���{�0ll�}ۅnJ����� �Z`����>Oy�hX���
��9��x��� �Ő?��Y�ПDM��)��N���u�"��ߩw�fs�C�������[�wMD�4�6��u�c�m�t�������F��VC��шա_�B�Iwl-O86mH4�P6@������~���<��@�3�g�k0�ϒї"!�E����y7����M��d`Z�
� =�`;>����~�h��Z�y�Cy��;.�����C�MKY�(X��X�m�x?�I}+��U>�sg�$��c
����E��7���*I�+e#���Ih�?��TS.I��eXӒ'���Ⴝ�Լ����%�H#��Q�+>�n͒����s4D�߳�;���>��z���B�s՛p]�!���c����`b�Ӵ�-(ə���NJ�Da�H(�[�~�#�(483�Цw�x`6<S(���_�fR)��˔�Jg�uZ���c��#Ƙp]�(p��^�c"Hg��Ͳ��QX�%���A���e��N~Д�Z��_a���N��_�&�0�ٵ�B)��1w'r�{s9#`�s���o�i��x����a���ӏ��	�$ob(7�W�a��_�:�v�u�w��;wI�_���,EKOmJ��p"��V��Ο� ����6?=�.�C#]^Xi�-̨�[w�</h�RD�N΍���`�;h���=N��b�s���S�4�#�!���u��U=4'�?�hMid�Nv����Mj}J,r��_#��t�l�f���6��_Ǔ)Pɕ�h��U2��ڢ.���@|DQ�w~0^_��4j���)C@,�.�+�Ȥߤ���襳��U91A.�䲜ё|�P�ʟF*�X�����}����o��	b�޴Y�O���uA�G� G��]�J��<��o�JD'u0���#[��r�h�3�XÜǃ=<Z�l�{�K<m±	���-��]"��No�Q�6^�Ow���c�6�s���a�e�Ճl@q��ﻆ��I��I�;�N�:j���g�_�pd#���~���?IZ�:�A�s�Kh+����BoÔ��*(�����e�@�v�N�Gf@Lx���/X���r�=�KR*�*��&��O觘�_7W6dqXҿ�%���X��W6�au4Eu'c�H�6c��*l�ؿ�|"���#��d��Q���e_G˷M�X��c`�af��ĝ9��:��q�
HQ��^� ��(��؇��pzq�r�I�0�iÊ$�=$Ш4C$ӑ ^��Rj�Xe�n9�X��KD�mN���p7��}P���eF5�����������wѳ���ۀ��rÔ6�ʀ�11���A�lh�U(ک����2$�IK�����	[E �-�!91(�)pQB��J048Ҽ��Ă�Gt��g��
)�rms!�Zf�2�LȚ�DbEFi�V|�,z%t[�U�!�����Җ�4 �Tw��gM�`Qҏ�ZA���|��O�x,|���c�+@@d����RN�ġ���:>�́�g��)����7�ͪ>�v)�P���*f(Dϟ&��gKX��Wҭ1����&/��u��3T�-�tyo��9�Ѝ������]�A�]�\�=��?�
>W��B�`0��\���l�ڧ����$��k��/�~������"d����nz
�%�S�R���y~v��Z��g����]���tj�$�s�@J'D�{�)">�@�٭w\<s�/�+}^��7HSO#���񪌁���=}�E�P{�ER�R5�� ���Մ�;���8l�sS'9V��	�u��عE3q�dy� �f�L��E���xKN�\w�/�3���Ov*�!S�z���=}���7�z��i'�FP��*��b���H[�n�ʒ��jixP(nͷ^@*t�8��r���гndƽY�� ���U����]O7�!�V0ǐ��~A�Z���w��k=�ћ6}��K��*���L4���w�˩t��7�ĖQT����Yv��3�cf���M���H�k
���N~�����L�V�Lu�����1WI�93�}�w����cq\��.�S�T
��>�J1�S�ƥ��m���Q�8�1��H�������{�<�,چ�.���.�ց<$�l�Y���^j���t�.�TU��6��F"��!w�N��xW'v��x8�^w��o�w�)b�#]����\�K��,�M�����S���(x)�M|��+ ����5���ۆ��2l|y|�n��8��*�G{�"%'��.t�x5�/���DOH����;XTD�|��e����S������/��%��|M3*f%ܺ�p��j3ml����&4wh 
��@�JO���'�����9�) ������֍6`!�L�n�m=��(�Vn�iZ��aԒ�]�7:�'�����"�p���l1����N��l9��i�K��ͧ[O��tҫ����[������I����Q7�y�}JW�9��)�j�*9�0<���H��dpx�P�-�-�/��Jܱ�����iBk��5#��#�S�Q5��Q�9$|��y�G�ɰ/�aj˽�}J�����޷X�0]۹W��o@�Ԋn��e�ܥdh�ꅟɄ8(=���Q� uV��ğ-g��l�ŠB����@=���/Ѝ̍Mx:���s|���	]�ȧ�n�XS,]gX��^l�o<���|6�� ���st*'J�um漠����(8�+~c �'-�hä��T�QA��zK�?WW�4����v��d��c�
�;��%�Zif=u�S I��K���	�ɐH�8ۻ��7|��n4	���)Aj96�� �A��j�A�D�{�6�L҅7��/(��u�}�seN�=�c�D��4"��� ��P�h���a�WCd��/I�]�ݟW��f����,��}�?U[��~��qs,���պ��D���rr��a�*m��t'���Pw�|�a�42�;ˆP���K/l�V�_ �}��Ϯ><yW��R�!�b4%Q�N������=<�h��[���X��R#yI�� ���1��N\|�j�A��i��;Z��]��'���-���P&��\a(�d���j5�k@gs�[y�zpQ���x�:�K
�y��(G�L�=2��9�)����4NC�+�Q�6_�2�e��
-��3,��T0�$hV���d�U"�9�b$.����ڇ;��q���鯵�c��� ��⛊l���/D���+B�ܓ��?��c̐���˼.u,-�G{�<nbPQO"����r(Y�S����sY �)�lG��4�Q�D��m�m����!@��K��$��wWJ��I;V�D�G�����J蕯�����
��f��a�ť��m��|�f��2#I��"/_��ю"'��x�:eM���;���=�SC�3�ā0&lK��c��M$�/��B�Ě�KfJsME�e&0F(T�vuԾ�N_�ͧ���I~�S;�n9�,;!b�ˠ!�#Re
�{��)y��QN��'>�D3JQ?���F;�`���-n�|���CV�} �B|k�s���Qo�G�i�_�OH��;��tv�}܇�F������;��88[�#l�;x����NO!t����f�0-��b�O���5�з������������ᜒ����T���V*�DBCo�� Q��4[w/er����� �k���<��=/��ɂ&��#w�̻�M+U�)+PO��#bdql�԰s����UUVj��ɛ�m�R�#�(����D���,�}��ԓ�R�͔8�Lw�`�*��_�QL�@�5��ҋ6����80�V��wp�b,$�4 *e�	��b0}:]��n}A̋�T�U����F�X�����&����<�i�N���"�ä�.����Kd#�����$�}O�V&�X%��IB�z~��N�ߤ����ߢZϲ�:��}���X�}I@��凊ʱ��}��dn�Q��d.�6&��GɌ�8@�Z;�{�}�ܸ����i��^}�j��GX�숼�x��9
_�LL���VOǟj����V7 ȕ��IV^l��;�D6���J���L�r�8��5�7�ф�n��)<b
�O^M����%]c�U'Y�$5��*'�O����En�*@���V�h541}�I�.*N�("%�Ǧ�Ndb��ݺ��Dd�6���z/��H�N�N�?���6�����ɛ�PW�j4<d��@��7�y*A��ښ��o�!�ٕ{\�4'b�Err��$NS�ʛ+��͜��[�]e��d$�>a��~݃'>���IF˅��BW���*�<��I0c��f��Iߝ��A7y���PdEӰ'x�Mw�R��/<L��򸮮Q�6b��\}+U�%p�ܝ�(�a��ަ8�����=�դoq2���(jv�&Z�;n-b����1����W�k뱹�u�%�d�k�{��9k A�rBKr�#lX��]>���=l�'���]�ܒCh�׭m����t,��@P!�)q��^$����6�(O�샕m�}"����I����<�ٓBu��� �����̲,��e��Jc�򸨤q@�T��D^>Dɚ��o9�
{k�����y��mI�*���Y����a��<f"�
����\����:�N��7j.������-����B����l7V_5���2	׌�����X���(b���C~�$�-����G�'���hp�$��x�m�kZ Ɯ��[W���P���M>l�-3�ײp
 I-���?0m��	⸾�j �Ml���ٰ��b+�1򛼤�^4�����6��y��"T������h�R�rF�<F9�s~=]]e�:-ZZ��j��$������~����S~d���P�S�⭑e���pJ�3���J8sm�L�u��{tTp�f�9�N�(}k�#"��4���0��[HdA��Rl�:�<$�Ϳۋhs�v�L^�dG���.������	��G�0�tQ>�Gp{�ě��,��E9�p�(�Y!��7��y<L�X�9�\^�o2�ڠ�R#�!��=��Xd`-�`� ���c��o'�ko�p����걈�or4lf�	�<(�W [�V��ʔ��B�9�<�8�JO�2���^�D�j,d](+��MV(�,�JS��Mt��s���rN�
���0��{]�>o+%"+��I?�3��E�g����VW��cخ�� %7,.�I��@o�iiw�Wi�?�ֈ�%���y'oߟ���p%���� ����?�1��بg�r2�߫t���X�$IV��zf�H�v��4��̾�d��Ԋ��[\��6�{�jZTmh�XD4�'/+焾`��^#S�Z�Ռ�UA	ν��ME�`P�Zsڙ�T�|/����*E������s�d.�'[@.`��<�WYZ^7-|��BZ�:�����ޜ�	m�4��#3�y���x�dP�``~�P ^]�>�7�ХU���J�7�|1���D0b�F鰜��v��><lg�+��t{,�p;Rzp'+���	ތ�"j�W�}� ���`^A����L^��
�Z,����:�$��@G�-~Q`������φl�깾�S��G�9�U�1�q�m�mPI��z��[^mnBQ�#=_n�·���i��ϙE$��f�e�����09�uM�v�R]�z�8� �����s�0^�_Sϻ�3_��<�񝡕WD�+E�`)�4D�� �%��8�m�d��ԳJ�|hp��iVOl�&�W��I��31%�]$6`Y��lw��[���/7k
���G�W����C�V�Nb�;��#��;�ɡ�Ӥ[�g�C�����zf/V����q�͘����`C~�B"�]��&=΃�ո�8��Q#Ҁ��i��d�3X��K�j���`��[�7�2����A�a��SQ=��ci�>|q�������̸dB�԰<�,���Ro��jq�ԗ�a���;��}썮~�_��Ivj�(>3�+X/Xoѝ&��q� /yG�S�c���Ȱ���y'仃�G�a��@2k�Y)t��,�U��D�s�t�@�!M"�0�����I�[$� b"-Q�Ԧ�I�F�Q�
M�wp�|Ȕ��� ���~�xԕ��z���v��
v�"�O�F��}����5�@\(�s������"��Tm��׬��U�/	>�A��+���rc�!\������#�0��ϴ�񝾘<kaYk�ճ'�@-#�g�=��m�r`UR���+U���Ta�Gx�Bx��|�!���c2��j�܈b��F�����"�b�0�([�U�3����[��^s`d���#e�Z�l����1���v��!).�(��{T1 ��ع���N$���K����e�Y�F���[�[e��`�D���Zl߱7Y����V�	�ɛ>I��^�Iw����j�Z[����!��V��h��7�ٶ���j�75@uJ�]��^�2�5��Db�,5���?H���f���!���WmPmEe�&�>侥$(mr���_-b�B�=P��0��b�Q�V!l�K�� ��|YCka ����:oi��$��,y =��(��n��Ɯ�`�Q ���@�!�7�0lUW��Ӧ�JSa�(o��фG!}	�>K�8zm�^K`k�<C2D1!�M}L�~���y�ir�S`�)ja��Q*�g[���%�y-��	Wb���ֆ�k���,�h�M%����w�5)��S�'���S��	�����˜���yǝ_�C��$��7#���T�f�ܥxP�&�3&�������ɾzj��c�v MYpqH~�7�BO5�d���PC��T
Ƙ���xf��j�%�A�&��&	:��lQ����ܢ�����[�%z�G$�K�Ej��7����6��,����w宷ڬ�����	�\����K�I�՝Ϲt�O9m۫+#�V��ޮ��J����m[{�PQ@@�j�?�w��"8�Ҹ�]����� �=e�9(j:��'�T�Z�����R!����7Rr�q�˿�<��eK�d�9��Y8�7������.x��J?,�U0���g�?z�9��x�����}�ؿU]�u�\��(��gnAݑA�@�<V#A���-�4�Jk40���v�gtda�;�e4�.�V�s>�G�rm�*��u,{T
�5��X/��B�&'\���*��Q���t����=�8�H~b��J�Եg�W`]3�o�o�O����ꆩ�G�e�Uu��C	���%i����MC�f�b�N@ܟ���3�g�#�c~w���ci�[~a&��65���9�����7�nܽE�?����1VO��C���3B�w�D*��d�2��h�����Zx����Hs�n|�:���K�+�B��l}�(�*�}Ʊ����18���m���{�%��"7J|W<>��o���Hgu|�$�n<=�/篗��|�Z�J�Q$`��A����8��^G���4;�)-�
93��cBmP�yFR���`<'�<KH�ȁ�)8�$}�f "��6��S�����C�á��ů�bN�^����0���'.q$ J۹�/�6�;q)�${պ����r�!�ik�lL���[��0}� �#�g?��{7h��;HCJrE]��U�S���Dy�h]��$���?a���D2Z ґ��415ˌ�s��i�E���ʦ���/�'T�ԍ����7 ��R�C�};�:�}<{.�����j�bl�]f	k�wӢN����	|gR6���m�;�[ٰ�:���$����������W��R�1/��[�5� �*�әA��t�u��`d���x2�7��g��H��arr�&տd�^��{ǲ���`k�(bo�;�A>k������p���1'*�
׼3
%��X1b�����^���zu�>CDA"�:b�|Br�lXXlxVHYEB    fa00    1340i������_(�M�����G��1�_{���YN*�pΏ}�_����5��?'���Z�O��ӭ��7d��k���Zu�ޓ%D*�m�9�������\����j�i&@GrN����$������0
˱4H�_[iԢ~�~�JG�,��b��4��Uk�Ũ��Pw��b�7\+��E�Ǵ��k1�)����n��Wa����.Z��E�J�&�'�3��8b �i"����1��_�8<)��Q�ӝz�"ӂʅ�����_	<���w��BR48_B�t��6'�e��������8���j{�x����F��W�H��P]
�=����J�=�t��^ýL����*����Fa��z��fw�p�9}��bd��hM)l��W���#lX����*��؁�g��r�Q�aM#4�<�6�y�)~,�ǭ�&:��Lcp}��D0TR�l���Ȗ���c�� s�K(&R�N�1	��:���jD�$�4.��g�'�ɗ��<����^,�b�%{x�m5�%��*����P�)�����Z��C���>������w>��.+P��*g1�Q��z� 9�8�
N�-!)=�W�`�ޑ�&�g5����K��VQu�$j��n?VREOӝ��C�_#����ڗ��"p��-2a-M�/�d�[GR0oP��A��Vfn��g�A�P�S�g��R��[=H�r���@�p���MRN���}���XKv��1y����G:P�����Cg4��>�%bx�2��^�7����/2G��̰�5�0)>�� ����A���.�?E�K���K`����sB�ߢ	���B�n{A1��l:� 
,����+�#�z���`����)4CH4`(�Cщ�K�#Z(s�/�wfvo��8�֝�������(��L���������#�߻ǡLA̡謱mL�[��l�_Af'�},L�h3�`�0���5��l�%�-�v�����T�z��
g���u��� ��c�;y]L�^(<&l���[����⇢G>�7��6��=���Jr]&r�7o�bJ�wqi.�������:?�vz�6��`�V��Iq�8�5��e�V�OTCo=xM�u�rWRi15X���q�Z���M3��Ș��,G,*g�ݼ��E(���ꉲ��[b��h���d@�%̅�c�Y�����C��ѹ�b�eH:�)���֞����`��C_"��ͦ(u��&��v>,꺝N������2��6�5R��֯����+�^A�l���3�b�)�_�1�R��yز#�׊��e�:�
��!(9G�̃�<3J4n��Oƕp���C��̑��^�ˈ$��j�6�)ϻ�v��:ϐ��Wـ�Q�n�$��5�Sg*>rZ����wk�D���!����;�'A�v�$$�}�{�t�Nfῧ���q�E!)��M�:~"G�?�������I�	|�}����̱Px�c�a���F�uNr?.nњL۱X�ɩ^BA�O�o���Y��x���)S����6��eQPB|�V�X��o�`���/�[����p�vTv�az�JEG	ì<	{����X�a�>/�iu�ִ.��SxЄ�\{��K�h2g��\�U��D
�f��*�b�o��a0�E����B���{0*�Εޤ�
���<±��W����^X='nb�@��;��Tp"�-�����Ǳ�_C�P"��v�3�sM�&���:�_tr�B�����a��OHk�#�\�zN�G��;�p�rW�lX�<m�ܞ�� [Y��sn'�ڌ� B���i�ydj��XX;�57h�%�'M��I>��T[�2l��� ���~��騸���8�ʃF�0ݞ�77���X�_78)�*1���o�%��Y`s�:�D�Q�-?2��cI�I�ת�Dx3p~7��	e�>ɏ/�\�|�]!Nَ/u�,����e���r�ؖ���r����( ~s#���Fb~l��U�UQVc����96qsX ��W�����R.xU�F"�;>N��n����jzl.�Lt�����n��cj�i�P95bK��g��Q�����>(a�l"�(����D�Ɣ5
�XP���d�R��mB3Y����i��ګ�?I9r,m'\��(3�7O�|ն�!�k�{{0�.���M3gr��y	+����A]���:�ķ�fY��V&�A;��
ۻC�k��ZD5<M�Yq����-�����`�T�/d�P�����v�����N8�=,U��݉9@c�U�f��M�U0�@�!c+q?����N^TE�5*vV��&���vk�@���ȋ��^�m�3����À��q�J(ɾ'���No��l�����&B�W�Lu��ۂ_.��A�tp�{���,(�A$@��5[��s���g����`ەDZ�eYS^Ap� �g��sj�M_1聰~&�Ɨ��qQ��x&$�X/���+��e�@!�
�NQ�����:D��%d'f��1�=XQ����C��7��tJD�A�.`���+�x'��&���;����w]�F����~����!��뜨1�\x�����(���(L�Z�C��%��h�Gswt��z2W ��o�J���#P�E��`��D\���(6ǭ��'�4�����x|Uum��{lߕQ �n5Vw��P	\�d!����d�Y,l��C�}Pj�{�Q�%�t��AD�^:A�h�ax��l���'hW��h���͝�&��Ph�;Q��-��i�� ���`86@�N��xe�P~)�ӬD�{��L�^�Ҹ���%�D�����0���R�j������(�o�?�[8���t�ՙ<YC�]�d[v��7'���ٚ���L���Q��D��}��`�`-��� L�*��͓���U��g$��(��\���I��+�"i[�-$�6=r���WSHumeJ8E8X����L���fo;�Ǚ�����0_�|���x�-����5oS�]w;�s$L1ɑّ~s��L@�����V	#¨A�T��G�A������`aT�^��|����kz����h�c�dL2��+��C�MWH<|�Ԅ3�c�7���� S�7�V�U�g��(�0��@���[��$ �0��S-ў�������Z��Ʈ5�.��Ǹ� ׅ��
1Ǘ�E�L��T^l�R���T�34�b��y�8!7]�n�e�v�o �O�B|��%�>4j$fw������z�}��d�Py��=����Z5_�ϸ��.jܬK5'ÐS��hR7N}u���w��0��3�P*�Av�xx��d�D���,5���	���%��MM�W�U�Z�O�e��-{�!���&���_qU�KL\y����)P���i�w�ݡv���o�Ԏ���(u�
Pr
si�<�'̘��|/�r }���g���|!!{j�"/�$�i�sh<��V�(���3���d�6dϰ6�q7�Cj�H�o����L+�c��~�D�2�[�O�s'`��c�z��D���C��&3��q"�e�u�0�p��i��^T��Q�`TN-�og����Hwr1�9R���$?\����/�P�*�����7���V'��c�E�5>	K�e��sp�ں�z7
���ʌf\�y�h���+��!�� 8�����)�p�.@u����:���T�u�.�Q;����aB�������M��˰�f������c��� YS�"����v�����~���/���G��Ңa$.(O<�9�y	���0�TW䗔4{>t{u�
�}�����/�x�$3H#K^2�i�1�Ց���!t0.=�I�<i���8Ϧ��W����r�&6x�P/�a��Oܠ�)ݸ��Dً�.\?�PcËw!���!�������j���=�&��Ey�)w���la��䟁��:��1^xA���k	�Y*j��u��2�a۫=� RN�e?g�i�ҟ}�5��.�ؑ�	R^�:/�x�^�:[�L4å�J���p�����r�Yb����xX|M��+-Ď�I8�����!�))��8 ��t&�Eƭ�̼���/��=!quI^(Q^!��>rJ{��*lg���fe|t^ކ�%�gC���݁'-	��W�pG�c>�H꙼Z'j�z�p��f	�K�N��k9�a�p������>�_�BL�1�QfO�i:�Y�Hn�&��j4h(j[�}��O+�w׎�I� ��� �,	Z>-~͌l7ʃ�}��JrW���w�2ə{��L�4Σ���'�o��죣7օ��ۀ������y`QF���������]�Ir� ���r�E��1�s�N���\3��z�S��Ў�!v;�[S_Re�ֶ���L���Dsi��T�rK�ſf!�Og��\8%x��I���p�K1��7r��f��j�u��&�zx�"��q�Z�1�K�2#)D�0��U�m�����B*o������9Z6`|������P��K�m3�O#4g�����R��˘�f]��n.� o:��b-9r���1�:��0�	�Z�����d�0I�C�MS_��.�L �Qq��^��A�❵��6-xk�mi��HX��74���?�\��Yq���E b+��0�D�B�q�#:��ϵ�d��N����ޒL�)'��HWq�H�NUA����������5�y�����z{�Y鉵=�@z�����w\�����:X�]��{��pU�D8�!�7�@(k���N��+�I�?֪�o����?[e���B$�mZ�I>�윢�Qh���0~E�殷�������\6D�K��N����+��Q�I��7cuj\�:djآ���c�xk3Z2��8���}��]B�q��夆�Q��<XlxVHYEB      e7      a0N�ܥO��s�ܡ(�/?v�t��N�r`<" ��d�״hZr���c�gޕ M�!v��������p����P箱m5�)�u,d���$۵�_�7!8;N�}�-|�/�m��̱i�s@����d��˪�����T�ԏ�%�?a�����D@���4