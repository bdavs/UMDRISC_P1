XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?L>Lq���	��1���y���Z֬V5Q�P�hF��3�M�ZS"_[v�;��Ҳ 4��T��< o����e���>���7���o~Ǟ��h���!�`��^~��,���`��.��8����;��v��uIQ�ГE��x�q빝���� l�y�O
�Һ��3�+�� j����>֬�mWs�pD�["Ѩr1{�J�I���wk%���s�p�ܯ������0jP��a	��zvъso�Y��m�����"m,�e�Bq��<�>$9�Dd�Υa��>:�̵5�?���<>f�<�'�PS�����F��hI���R�4�s>�1ƾ�c�߂�������䞒�˚J�>zR@�E�Ā D�y`҃�\+\NJΣ�q:.�%�ٟ�-O���Rdvr�'�ۤ�m���*0Kև	���u�/`��o�����@2`�gB!["Z���:Wq֛R�,��_�3�E3�C��� ��]'�A.�����F���t.l:ɗ���[h�����f������x-�;L��%ǹa�Lb�<�	�DV����o�2�CX��o�%�m&ۚ�A�T��^�D�d�k8|��P���$ �q��+���!'��ϟn�[����\/ـ��C�d���Ŗo4{�1b���X�Mr��Z3�C�|��'��!��3*��)T�+w,�*�"T$u�נ[<͊^$�j�!��ڜRW� �<��i��Y������]6� +/XlxVHYEB    fa00    1f80������p]B|z��=.��yb9Z<�]N���^�6��,q�e]��qUuճ�.,x!��*��g��P��do�0c'
Ǩ�A���r/`��[1RLX{I���C����%��b�׻�[.�_aH�T�L%K-K׉��Mǁ�*y��@ב��T ���������nJT.zv����J�67�����$B�� ^��H��:{��v
C�Id�ds��6ܬ	����pO�!lxs*`�Z� 8���X��6��<��4�|�I�Y���@?г��5	W��G�䨁�������
�
=�Op��kX��0;��	�)���u:�UdXU�yw@6�a��T��׉qr���5ԁ��5e�F9Qa���<&S�y��M6�`�N{ο��#�����n��Q.�;��!Sx�0��4{j���1O\�<JLZ_��l��/5��o��ћ������
����߂x�e�a�$
徰z��, t¤A2�U�9��< ��h���h��ע1���󗙃q����͏LJN\��#Вa)��DH��Wll�TFϒEӿ�AE�0�A��:Pn�ˇ���)�E�bΤ٥���U@2�N�uc�xs��s@�������d��`�Ρn��o:/�J�1H�O�C�b:c>�i�TЎ[~\�v�\7��_�9t9"�f�"�uK2�&z����2v8�
����CR�Q��sx[����S�� ���ۋ����f.�Z��"l��1�y.�`��z�>��!����q9�{�cJ�Z\H�@,ZX�m��G�q����1�{�z�>��8i��qћ���0M��h�z�,,�w�]�30_�!y���E����S���P��Ё�q�����.�E�������"T�G-9�c`=;�B�kFlx�@j�7�DC{�m�c�3��3��P���y�y�G��*�Af��QG�5�;��
�A*<Z&RR7��B��+Q���p�'�W8�vEX�+���[4a9��#!����tl�v��Ļ�-��,3�}�8J/Q^�F��Z���3��Q��'[*���>"��^qů��r;�h��g��#�"�+�X6x�3@F�-
�j�=V���=`Zxs5�2�4;Ć͵���w�0G�9R���}Eѹ)��vD#��� ]��ڲn7���;��3�|rq����<��d�}U�T{��MO�	Ԙ=0wL����a���'�P'�P���SA����w#x���;��|d+����m%t!�q����u(4�
|���>u
޼��n��{'�p��+�s��R~��4�ѬF���銖�r�c�hJ��ݞJy�n%|B0��\������4�Ѓ-�{�RJ��	ϸ���ݾ���^̙�"�	��"�MLA��"�/��5̿;���Vw�3ؤ�|p��>�&�c�&R�6�=TF�t��6 ���h:<�^�VPؐ8�`�����"g���p/�F��ꠋ�*�$yմ88o0Ϗ�x��j}
<�Kky��,=)�1�� _ȓ�����L��-�������XP���k�Yn��ƛ���W��C���uf98! p~�vh�3�ѧ�~��Y%��
mb�����Ǵ�Y�Z����&D�/�.�&��8���6���56�G��n-�m������q�3"���7ݑ���Rd�!��2bb�h:	w��tU֦z��1n��z�ku�_����\�e�y��B�˴;E�#�|�^T>�8�[�k�oI�WUX���8�	����b�{u�\��&{�T�t�A��%T)��I�����v�����q���L:n�:߻�y5�tgL��Ĝ/�Ǹ���.;�����j%/>����ҔP��sHkK��(6�řΕUL`�ٯ��]PA�,�����)�ѵYý 0�X�2ڊ}߹v��Uj��סU�������Jl;�XW��J��
xn�Je���b���d4���#7V��F1�
��-��ͭ-�_
�>4*�c��"�X'�|'k�����"~=gJ�#ڐ�ӄ�Yc~��zI�	��$*�<�hy�c��M&��	�݈6{��v�ِG��5Æ�e|��s������7�N�O�S�o�7S�8��h9 AS��F_�Y2Ē���]�����<
(��E׍'
 �a�DU�cƣ����>��U�3B�>�gJ���ᾡ@r&{�Kwg7��%y��tʍ�
$�)a�����M��W6D�l�Z����<��-<S����9�	�����v��Gg���f��*��/�zk4����a�j� �P���;b��g�[�u�;�[EN�@�S�4�kؗ��!��!�� ����T�|�|�>b��\JP΀N=�DbD.<�(M�*N��g(��y��'Q?!��[Z�Z���W�nl�mnP�`�!�U%��`����qӡV��XQ��\��N�8�=%��3�?7�t��7yX��2�����O���էaPq7�� r��l�M �9���� �g��TtT�t<�7=��j�y�9$�"��c`��8h�#��+�`���
c[B �(�g�p6���G�%������=aB8�	v��?���31{����-ڐNH�k�+H.�1����E׍q��O�?��2���O�ӎz0������|D� �;gC^-��;�!�0Z���w�oiR��#��-=��,��ir�w4��<���B
�wL���l$��$)��8tB���C˻9�?�эa'��z7:y4���X]{a��j:(��J�zӃK��nĲ�>��ųa��Atk�L9�����>�y�4*����.%o�>�LB�"��TA��%[#�F�0�薪�3%����eת��g~���m�d�y�FK�'MY��xߓF6���D� C����_$�W�����[��q�Տ��I�����C�]�V������y�����?|�q���&�*O���[[�1��(�\j�G.Cf���٥6E��;㓣j/��fٺ�ob����_��v�J�\��	�e��K �>���^ˢ$��^�8s���p��TA9m�D���m�ȷ&[�ԯF}���w�b�-��&7�b�%�eG<w���rG�����z&�|M+x��T��4�i�026t%���U"�Z�̝��Y�� �z��Y���l��R2%�]0��'���T1�D��Bzm��Z��n�_',�-OVl��F�}����}�<���=��io�k����{'��[VEF�J�@ikB��d��=R���>���i\�����8bLC\����;Z	{� 㧍k9(p�|?ҡ�3�b�p��f��o��@��f[s����V,.R�V�ru���h1���/���]�>����K����
�K v�����3���y��Xܳ/��.�^m�"��� Y =
)���Mڿ���2�����h�=j��3;Y�N-*���XeV�V�-���ݙV�Մ}�+�]5�F���y�F/Q�C?��`Bj8z�6ǎ��;Y+H���w�@a�љ�r6f���e��7m�HÅT�f���4K��nx@��7�.g&�8�J}��������z���pR�F�=�z��D��a_�p���Mg���
�l��.g��Al�
1���Ut��N�\����qo�����ŗG��zV���ɗ.����oy2�����Ҩn���wݻ����
ϪډC��zָ����}tL�_�,{n,��1!�+��x1�x�
1��E&��l��pō��\�
:��j���^WkRmnZ�% ���܏.u��VJĠM$	� *�S'��	gi��x��l���U"7��V��Ѻ�D�z���[>k0��@zw9���̦AG��^R�K�;�t{{8�O�c #kNvR�a��#��Nz*�T�U��:
r��c��ᒵ:��f\ a5P����>sq_�TL9������{6cY����}+^Y�y���J�Ӊ���يu��{�y���ME���Y����|�vz�[���*'�&�4�	!����eҾ�ja�-)���r�p��җ� r�ŗ����
֔�K[$��R��) .�����.�Ĳ�, ���I�\}�:S�~'��p�3�Q-Y�4X]4e
�$��rP�w�N�|�G���jY�����`|q"��\�F�Gy������˹�AC���=����]�,e3��Gm$gW�zJ1�d�W*t�_��jg��]:Q��J����a ���D��*�^���G҃�d�2�Y�K���Z'���?R���w���˯��.����c��#�Qk���k�=��H��^0=)np��� ڐ�q��1}��7����KJ�w�;����ff����l�D�I�`�*�:��2�j�0��!U�Ǫ�W#��:��tbx����K?�u�q�@�����y���(6�E@⍝���̱@�,��E&��}�͟o��t�M�<��5C$;�� �4�Z 4
#��Js՛g�\%h;�%SD׬��.׺�F#,�IX��1��c�G2���{&[�Z��9�erJ�Px��ԟ���*����%בIH\ۗ��ȝ�)�_;�/5�EF���Z>@��dk��ӶϲG���� �jA'�i�32l��%�M�!�E����r�.J�Ȉ��[�����~��Q���2�u�$3�J=���m{*?:�*�/aD��ޱ��x��a ��ES:$��2�9��(�����@MYJ�0�ud{\/E��^��+S�8�[z	���(�&mn�k�V����6+�}K����<J�9A���·�d2R�v��%i��_�����?"(P�N�ǅJ-�tȚ���W�-*y���Xh�O4>4���j��r��:��.�:X"�,�c_@�\����M���v�p�v0QK_��%���{�HQ��A�,8��I�T������ʛ���o��Δ@GB,���d��X��u\6MфG&w�~��.��Rt�A�n��Q�:�k ¼C�H��0C��#6���C$e������C�S�U�ݍ�БፐK.G	>Ѣ3;�%"cR��6o�����j+^�h���4���#���g�)w���6腮JNE@WL6JO�pFH���)��Y�����3g�qk�d�`�e8����&F�����|U���*�W�QZ��h�� Q����1V�'����'u�3C��2PH�ǟW|3���q��Z4��c{@fV��1�^W_HQ��7��4���du}�SM[&"���m�st0\�Bse׿���h���VRZ�yER��8y�_a���c��R����J�Ċ���c��!�h���2�f�&�EDQ��;�f,��s�O�LQ|\�.:����@^�w�l����S��1��_��Q�� Gq�6��3�p��M�YjH:	��w���~�Gp�� Ei�;�������9P)��N&.E�������{2�@yej'-������n3QE��!mr I��dF̋�QA�h~�&��E֌�O��I Qi�R^l��<���.�Rc߆(��ǈͰr��s����B��a�l7�����Izf[(�\D��9���4�݀��N��
��R�>�#C�;IA::��6N�C>L7����~Q�]=o������ʜ�=��WV�	B'G�O�����>W���R]n�4�w��4�w<�5n��''�DX�6E���,sk懓�it��H!��dqjA�vkv���_�웷s����n��3��N�&v�����c7�8�L1�Ӵ��`N��7�N���0ռ-ґ:D��N3LO�W�Sb��}��{gby�3[}�,V���W��Z�s!�hT���{���|\&��zp�`���I���C�=��*֟�5��R=a��T�k����{[���IdR��INaT��œ��FH�S��_ ����p!���$�l2�sc��D�2�`787e��n߰��s!"��g�ˌ�1d~�FRB��&~��܉tҝ�D��d���9����rq�yP%�e3��ӧ� n���?!Jgk�l������
���c�YB�)��{��7S.rJ�r�@l����Oy�C�3P�[x�6I�`��	�k��b����M`�P���<�N[�⼶'�fj��Jla�<:u�?,!|@(�����E�+f��]�r�Ē�*�����=��;D`Ph�r�R��=u��_C6{f��ev��h���dFc��#��y{�r��X��4����g�іEwO����?�*٣*�)�Rw^[��~�[W�����ϠhM/���-<*�y����E4�;Z�g�i\c�n��&���aE�so�%�Q�g]a%*�1Y���I�=n�S�>�0���&�h�U����ei�L��?g#B��hא�ns�cr۠��t#4k*g�� -}s(>�m�I���ԁ���l��o�{��P��u)��� %A�.������m����4�س�P��v��c��C.Pe`��a�'�Z:+�G����%��8m�v	@�lE�9=?�u�8��!�s��L�������)� �s��uP�=j������E]�I�*�X�����p1I��O��ÓӤk���r�3��#[��۬��ynj1�27X�95�V$����5�\ �}��v���0s�T�����K���z:
G@Ʉ|�y�[m�x ]��w�s�{<�4M�b�6d�P�$}�'��|~Ty�I�2��(6�8��2��C��?��z1[�*��a�ɧ��qƛ�u�"ʐh�3��K�:�X���d��`��YDb�k"���uN]�o�T?P�٬㩎Q��	$��	1 ��zE�u���]������ I��p�v�s��_Tk�D��%)v���%T�����h��@��A�K�S�,a�@����Uo�m?e��������N���YP_W��Jk#-�%���T�_`)<l=���?�kڀu&
ƂԄn���0����) ���#����ȼŎo^4ȏΐ���li�d�ݛ@K��ҩ��p��~�1����X9q6lt��%[J�����.��m=���\ޝ��Ɣ^[��^��S�V>�<w|">�Jͦu���+���[�m��� !)���?!N�ʗ70��ZwA�x�V][ �*o�Ev"�q= �s�\m5�W���p��pd�Zf�Xf=��ө�R�VKTX ������e��2 ɒ�*&��9-DH�I+!��������N��=ı^F��(8��p�I[��t�2K�=�`D��`ĉ#�T7D�����}��=�FQ��n7�VU�)�,n�2��g��ǌ��*i�����H�������_pY{���׾�ks x@���Ъn�s)E&�!�,}g���Y���'/W���m�C������m\R�L)�t��ޛ��~;��M�'�B֗���<���)��]�8L����)��8׉g���ƒ�E�'�b�S��-l���d�[G�7[��î�e�G�tV�:zMyQ@�j�����~U��od��^�]��b��Y�P�
�0���^�Ű����'f���$-����;w��ߴp1*�L�����9G��`5M�
�-�r��-��=�
ɨ[|�N��)&�G�pY/ְ�C^�s�'>��A����\N��@�c��k'�v)o'�e6�����%���Ia�aqMT]��N�-��մU_��Eݑس��5z�c��(������.���Z����U�?Ė<f�1;'oX!�
UCѱ�@����iO�e�6� k3��m37aM%IY]���u%8% �c���}��)Z_	�b=�[�cf7Z�0rE���r�*�!߯��!��d�R����t�ps�+����#cv
�ޙ<���&	N7��W_sp�f�WC9�����!�:�5��Jr���T���`�n�p7�_�B?��$����\߇1#��oV��Z��}c��n�3�r����HXlxVHYEB    fa00    10c00ex�)ǒ䃂\=#'v�A|c�n�#��K@}4�{~F��,��"�	^2�
-�2� WmmV�a�ג��5MU�1ֈ��� Jo��1>3T�Q��=	& <���\Eu���������v�T�B�=�&��S��16�����|P���_���8��v(�����_�B��Ȱ��	0���|C�/�J�E%ulԽ����B��S�(M%΅<���K�ND{TI[5ԇ��(�v.�a�Y�4	��Z[yH��0��A�c��t �M��|�M���,���b�X�lJ�M��|��mО$��W�X��ʙ���j��́�;`�f�.2���M�k�!��(�lў�Πn7���-k��w0t�����"���w�fl���g���N���a]%�>���T�I���6��X�
w�����oɛ�h��GaEA��:�ю��a�+���'�h:P	d�Ű3Cɡ�t��ߩ>����!X����Id�y ��I���֐��(V _夕�]�=V4��P���\ �CZj�=S�Lc��
�Ǹ�7�ɔS]Fm]�� ��J�=�g�BF�}�ѸY�qd,�5?NL_�6��>�8ݜ{G��¼� Uwm��μ�-��Zn�6�E��r
f، ��-)���3��N���8����ջ����$��jo���II{��K�a�sB�d=��e4C��0�3*}����f>N���1�V�Ɍj�Ñk�{/��fD1������)x;7�}=$mۗ?(dwE8��9o|yMI栛�����]@��k��~�t��J��N���\�Z����t]Yu�d��_0 ���^*�?=�@l �WW"�8C�vX�[(����z�	�ÅџW��	���X���\�u{ҧ���8�i�=*���Y;}#��c�0�%�;���KT�mU�p����\����T~jM�pR�>�V�_��D�/�?��y��-6����q����$�p[6X��Z��Xv��1&n>�d	4��ٗ�^����f��>G]�F�"�A,iCͼN)��3d4t2Ws��<\�A�Xܒ6����2ߙs)���hW�yX�� ��O��xO�8�; ?0�n�t�*;�U�?Y�u$�8���R��d3HWg� F&��%x-A��VU�A�aF�a���	�o��R5�G�mkT�7u�4T@	h�LX�@U$\��:�)�83F��F&���
\&�����N��;ǘ���?��6�o���ܣe�thB�W��	���s�_!���U�D5Ħ�A�d�ށ'6򨴶����U*�6tA�[�-���)??����?	����N]h`_��V�]�8���uCcZx �ݛ3�O�i8@��D�9��	��A9s�M�dZ� ��9E)y���8�3�s!�fU�I��(	�P����ME�/3p,�`1PU����Z_���b��[h���QD;���j�����w�l�/ Y��W>z���u�*���Ǚ�O5}{�����hQt����Ί�|�gÓ1���b��>j�9�xf�Wv�~���:���o�kZs��溒V�uǉ�����}��` f�͖@ĆK���E�E������s�׸E�`-'F�]��QB��;�T�� ;_�V��:5YQ#ԝ�9P`,�s�?QfNw�1at,s�p�XȓmW��o6��H��ǂ��r��Qye�FW�t*��e~�hǦ�?�b�L����[�´.��.`�^?0L�m�2�(9b�us��.�Tk}i��B�S���fmm6;+`��S���v�=C�|�Y6MvPB)q7��`ݥ$\v�(Z��~'kZ�-�j1M�2�a������2b����^������Y����v��5@CG��</��uy(YJ�?����G4\"���D ���S����tEC�K����+e�20N6����B�����:��î���Uve�d��Q����{s,#���L�-���#m>�m-���Ss���B�-Q��}t6��2�iP|��%p�ApČ�{�An$��*f���|S���}�=�rz��6�*+~���:4YNْ�Y7����C���x��E�};;JK���I�6bqoHo��\��v�o��q��m�2'=@��(��_�E�����`+	���F\��hǞ�Y�/�O�����k�<}g��%Lg�Ӡ�^�~Hl$��D���fw�b�����W��[,o��6�� <L�u�	��J��ˤ|�V/����������|Zkj��&V�5�?D���]�m~/*�
���@���������N��-34�����:�?E����?+��>đuKɨw3��u��r��q
#����m�e�E�aR�o����̌yN"�?O!K��#gU�v˄D�5����T�L�q�*2Q�ӿ&���{�nÁc_jH�<�r|��!�}�/8�n^=l��ه����OK�d�3H�!�d�d�:����_u���9�d}~U�����Y8j�V�ƮG���;^b��ꥦ3�.��y�#-��aX��*>M�u9� <�4�U��Ȱ�Cɽc5��׮ܠr0a���I�=t�tߺ�+���}_���K��!A�'�4	���&u���1�؜�]z�!i�gi%,�E�*U�
�g��cC���Ӄ4�TȆ	��`�����ސi��Pm;Pw��Y4�ǥ���yA�}N���٨�j��5>��:�/b��:���{NXVЄ�?x=_��J�~�����tgV �(姤�$#���/�����>�C���r�b�N��|��Nܾ�X�D�����8���6$�4�Sk�,�zf�t�΋�a�U��e@�d�s�2]Sn���j��0�L�B�?�l���e�Oa��<��������D���դ~���C�`��)wbpO�ΏO*�4��c���c1[�2�ɕ#��1�Q�'��^rO����p>�bW0m�?��;�A�fb�Ր9k���XV@@�b�ESF�f�ȵ�-|�*���e���_j��f�	��	:PAvF���ĞI�Ĺ���4/��\\�4=Ymh�5�����,����E�_,�$h�+q:��o�}���s#� /����u`�B��ԠBz.k�Q�Z_,�a�52m0/,�$���>�=3�pg/0���q�ɭj�R�ۇ�L�bu��/%|�~��&��������}E`�;�mL��Q�N��~�(�h�����	'�!Wv��Mg�)W׌�>�n��'5�v.C��@=�L�� ������9`d�j�F�<�RG���� &���&���	�TZd�͏���3i�Ba�h~�F�-t��nbo��)�o�hԐ)�݅��vO:P��Ňh���sIL�����/���h:HbK�H����aFL'�Җ�b�Թ�{y�q�k?X�� b��a�����4cC����QY/���V���%�l�(�7!:��A��.�s����{�h�YVv���Z)�TR�i�k�m	ߢP�2���L��.Ngr{����=m��5 �a���D��iM�e9���T9�d*��{�)��ЋRn�+�(�3�x�t�r��VG��ǭ�)Q�<d�Ѫ�E�	,�ˏ��q��p���o�ϖk�d����tUF$H���c����Wl��R~(3���������j�S�����8���qg�+�1�!0�¦!٬�0 ��T�m�fwVEʪ-Q��T���ٝ�=�=�Zf燕�Xݨ^�{�"x���Z�}HSP�O{P�QI��t Q���R�d��!��VEP^�6��@���e�SK��9ZG�"P�PS�~VJĽt�p�1,{�[_m74%�w����/��Ar%�2=���<��ĉ�Sq�߮�2o�ş/ >�M��u�+'<��uۑl�]T6Գ�k�?�_���:��;�!�w���S �#�7�
�bHyWJN4�����`^o�iۊ!��\ ������d�9��j��tz��H����f<��4��ڇ�:������!Z	�x�B�b59�!�__u�i�W%�&ָe>d�pn"?{�|ˌ�vR#���3�N�]���.��N�&��ٺ`0OV�o�5C�<�d���;�����$��؟����+���&����X�t������[we��qBy\��b�@7�O)�x:����F�X�c�Ձ�u�`O�G��:bM:j 1!z����=u��H�^��6�Ę���GJr:1o���F>Y��ϩq`�D<7��Z#�;J��>�l��	��<�R��4�n<BM!ňCl"0��@�V��g�c��XlxVHYEB    fa00    1140�S��;
v�ѐ�ӵ���>��-��:w�q��V :�@�ʗ��Կ���O ������k���p��(t
���oS��Fi/����)����4Ʋ [��|����M����E�i2���� H�Y��06k1�`�E���c_�C'�����~������xJ�4����\���~^Hn���^�O�������E��R;�㉿B�k!6�p�vz�p�?>(���G��u�$4�X�[bH>����qX���ϚFA�r�P�=2�q������Kb�;���LS%�㼙{_sl��S*$�b�5�@JLqmt����7YVo�����t#��E+�̩p=�K�F�.�l|C�3�y��x�����c����F��F�ǀ�}H���t ,o�A�/����)_��V�0<rY��|�J<�?e����cX��!�o�@C�a�0�Wv�Z�������2(��Ԟ���Go���<ɠ�B=_����W��~�(�O��J�g�飫/�ǅ�4�.���3��z��5�욠£�WH@�RHS<����G�(ף�,��2��9#��J�W���	cU4}B�D�e�?v�i�������id#�ǈ��Q?�Ǭ�-o������j*��W[7��4�Ɍ�E��q��:/��
��۶�#�[�jW��q�g'�t����;T��-lC��둚�\�Lɍ;PH�m]?ؓrq]�` ���)?95��� ��W����Z��Pف:�t�B����Y��$���g� ��U�g�W�z��l��E�M����r�fXLSd<�w!|���~�d%~�?�1�?0UH�O Zվ�3IuݴM�}��aKeC�Q4�q9v�h��;�R�l%������m\4��Vx��+i�
���!�긟�Oį����'��2���4�98�1�I��g�!1�%�{�m�ᐄ+�`b�;^������#�l,'b�#�i�y� ���N�5w��A��0�~���#��bhP��/���+58͡�A�DG��D�����~7�������z�TA��~C:��-K���_f���u[^� ��[�����.j�;%����b���Ґ��|�q����~� ��d�4a郏����XR ?TgG�b�u:	�|������8;я7y�p������]}�r���ӈ�_B[	3��,�P{mH�i�v���������=a�tυ!E���C3޹c?$��b�%�"P��[�%*���~r��M(Id)��=�/��'<�b,���l1*�e���q���m��M�(T�����#]�|\d��z�� -��)�6���λ-FIv�0	�p�C��>�T�o���ż�e[n=T� �qv����4f|y ���@��d��S�L!�	�eqǾ��<�x.O<�98�
v�&��H�1H�W��ķ��{�y l&H}3%�IQg��	5�Q��{�g�iҿw�ׂ*�~*�1٦�W��m#f%`;�+��t��5�|�1U��_𸒶�b�ۦ���|��A��,�D:]ܤ$��<d�;���8C/�x����*\)M%#8ZV	)[)v�잁���|�u��Z�^�l�D��] �/?�6�7�u�!Xb: @E{�#x��rZ�;<��5�1��j�e�k��n��R�S';�Y��I�\V�a�=,���'�� z����Jd�U��hé[ZZ���D~.���W�:���I�`�9�	�Y+��հ�O�Ӯz�o�p�g����� �)�:��Ӌ���O���	��?�=���N?� �F	.��A���V~�է��
��i�g��J�[s|�{j�|�v�<���rԥa�?2�I�h��-y��[��-	*5L|����	�]$e@0�e�i�s�Z��Ä�m(Z~��,��m�c�V%����e��m��@�j��l&��L	����[*˖�������.�G�ؔ�����϶�� �43�����*��]��T#k�������sh���EHNF�_*&b��,Ul�Edx�o�/c��1��pR�IZUs2A��A1�`{}y:r)]�%^P�����@��Ǜ����
P�]�*�aGʒ�i�vY�Nfht��m`M ���&tC��y�#�:�E2�Q�g�<鬧_��B�=�i�l&H�E/��l�AOȧ�����x9��������
����������#�M���ȡ��a�'C#��}O�&�}˙	mr&r��вce������o��k�xg'�lE0�l�,�R��ʎ�sa��[��S�x�l�s M�+�Pbɡ���R��׎2��G3%� G���-���yC2�����Fe�)m����~��t���ՠ��V3Ir%�>�����l+���O����S�� .��S�(������o��Uq�O�g��W�^_2m�h�󗶑�$EcV)e�����:��z$!�Ī��������,�c0���ՅӟqD���tu���6pr|����b��sJ�wq�;ށ�� \\	�<���d����dֿ�H�`�}�JUL�"� @CdP��WzP��~��#;��w� ]�`z-7��(���;<���W�΢�h�x(��HT�J��&�(����W�t�|xǺ���?E��%���, Ń��v�и�~��O��?S_���6.�����BQ�Z���;��?���]P�����@��2J퓜卄#J3��i�t*p6}�|Ʒ���G�J�JD���4�X�^����mh�M�Y:�d��L*,��Ӷ�*LV��E�@t�8"Ǆ?�E��=�&b.�%�h��N�/�Ɲ��î��|lw��ۚ|���#�@�%b����g"S�P�ƭ2�`Ǹoǽ�s�7�2;Bk��@�qk8^W՜�:05`Q8���`"�4w^(�+]�;�^l�E�@��7�S!�����-#�>eǯ>���Ҁ���t��^�4�P��1����Ֆ�E�Ufx������т�U��*.�Nb�x��r�Wb�Zz���_��:A�������Al��y��aX}����HnM��<�L�B���"� L�4�_�p���(�Gw�Y9�l����ʈv39�_�}yR$� ?+�ˡ{M;�_Rw7�.�nº葠��;c�T�j���2���kԒ�S��2;eu��XZ��b����KG�Ksw���]t�X�J��&�N+).�|#}�`xE(_S�D�ߴfvT{��Ct_Â��0�E�/�� p�Y�H�2�=�K4c�;������x|ŝ#wS��j6,o� I���F�g,9Ys����V�I�o��|������L�l�^��h'Qxߢ�1�|����C�[q7x��t��!�6R���7
����BTp�}���/��h�N �xv�w�I�/�7�{t�ՙ��12�����w�Xu�����!|�9���}���;��Z&k���*�`�������(��9��2HH�ݒ��|ʓ#���t����`ݫ�?�jb&+���8M^J=��FK�B$�q�������aҾ��?+F��s,�ٹ*�>M���$�5q��f���&�%S뷧|2i����U�o	b���P��Ȣx� $����M���t�'�v|�gy�c�c9��E%�b�\��R��08�@O�ٴue��6�P�/�_�=��7�n4]/:t+��#�Jy6W�Q�cy[!Y�lp랑#=�*��;��G���T��Þ�E1�����1Xb!��o������˻O�jJ+R�.��װ�w���F2��dᬶ2������"/�~scM�^v�:���Y��OL���5¸ gݏO�3ޱ쌣1�izʬ�MٰP�E�,��� KX��������tټժN
�2"O�����<�PTՌ"-"֡���T�TJ��IU�1�����\���lyH�޶K)}B~@�ε)ڢ�� ���.����ا�fB
?��Eql̶*~��� 'ƥ�*1z�'����T�0+[�	*��F��/k�;M�0��YD�����3�p��/	���r�h�a����v&;z�`K����|�!&�^aB�uq���Ƚ2�@��ҿu)�W)~L}���A����|�w��۟���0EMϽUr�G��9�e2�'�#f��0�F��L4���,U��SP;�!�fjĪs��e&��ij|{u�ȶ2���x��z�\�3�+�bX����Ff{=eY0�|�q#"P��1��Z�g�M���@�'� 鞫��V��4��Y��!hB,��lw��2Ϲ�/L�{�|�����,r#Y�ZJ�!�ʃ
�>�����G�1����ˠc�.0���(�.�)b�����q7Ћ����g>�É���ͽ�-���+I�^40���thEXlxVHYEB    fa00    12e0uxK�h2~EMa$Hy^�ŋ%����ґ��w��z]5�%�ufh�P�k��>k���<������P.t���:: 0﹁�9��\�{w6���b���|�%���9m�v�ҍ?��s�\��S�-$0�C��XVxh�o@�2�|�l�ka+�=J��%"oL��8ۇ';l�k��ۥ�!#N��4�$�nF�/����|�T?ru��^N�J�	D˦�K��Y�إ��� ^�p�D�����^pdW+&Q�B�A��(W*<SҚM|��W�^��>��2<<4����A��-�@�d���R���w�%�,�s^w�fA��Mi��6�a�4��3�VJ�y0z��QLG�dA�J������7X*)�ϧ6
���^ߐ�V�?
����ύ�_>�@;4�j�-|������kb�y7�"`�GtX��4�$����)�����K
�zi�4Z#;U��UkO�ʪw�)u�x���/�P�t+Fdv�^R�m^C&�'���D�S�9"�s�D�N:��5\m�����}�������??0��D����"���:G��q�����)�ŋ��|���܊O`��?���j"JJ�;�H<�&��|�x������r����'���3�T9w7C1W���);��9apx��@_E��J����ϖF�J�>�'�	H�67�?M����o0�bB�XMz��"�3}��RU�&e��X!S���7:c�T��}r�c�*?֚�i!��!
Fsa[�ގ����\�O �?���|�č@�_+�n��u�u�0W���i������Oxu��m~�T��
���ہ���]�z�i�L�]�@���ID�g�~�gя}��r� 9�$�yXr]��xՏ����/��6㖂�"�7=������+���$xDvpz�bc�WQ��̋����s�#��%F��Iz�n�Y���w3%G�A�Y�V2^QM���E�&m�Y���@�J`�|��Ğq&�z�~̉����s�� ��_t� 4OE�'yP�7��'�,�"Ӽx��.�
�,O�{�΃�O	�(�J�r���S�	�ɕ%��_���sTyQi{�=���B��i�d˜�zI3H��uT�ܬ�aZ�4�g��=?&cq>�'W]��7��;7��,��+p�:V��?iOu ���vY\��o���`�?8'��t�=��\�;4:�Ǜ��tg����2��ݓ��h����lq�Z��s�^:�Vz�M*�%:��-���ns�S����|�q��7�ҝcBN�U���2���l_k&����MMU����@W{������Ҿ���� �fE��� �����zE�c��K�p�<�����j�tw��T��L)�s[�*V]}��.����G1��FQ%�\�c�Q��ek&7����w�^ٙ�(�?:F�㼴���X�2�3�_��8N�&��.[�ۃP��|�5*��Pf������<Dm��HF���<�I�'u���>9��_�In�R��'#���MZ����4XP~)�G�|	��%�	z�yA���s1^0Le��f���m��B̵�`}��G.����-�I��8��e�In�ù΁a��.��߻��wDO#��y�CG���@���99�/�@�v;�??����E��%�i�����J�o�1��'n�n��H����R�6/��Ѽ�*�ӯ���;X��M_���}�/hY��A���<��\��|�d*A"HZ����e�},G��'�P������{���kψg�X?&�*��g�'��|e/��n�q�j$i<9':Sw՞/�{5�Tg��'�̬'`8�<"����VD���I��o��n6V�&Ci+��~��yA3���yB�V�R��VK�ef�-���}ʍ��<�Ւ��>XV��6����o�����F�ֵOXr���V�@:�櫞$3�o?h��~:B�����{B��V�c��n�O<�`�����b�Ý
w�M��ۥb�h�ێq���Ӹg)�>�.�5�ц��ıW��zw��'aV�����ul��j�
�|�دj�n�E�r+�%�:	.G�z�&����	���Zo��Y˭+3m���n⬝��6����/@�����n��M'���6�B�<�ֱ�-���U�A��Gd���雡6�i�i��57��ɺ}�L�?��e�����q���&4���V���U�P�(�-D��ڮ�_�&6+4��ދ}�lnBM��B���53M��[��G�:�W�95��`yG�����/�_�$�l��m�yQ���]��)�p?���>��ck�9��rc�׊bkFU��*k�X@�_T��פ<x����B#g��uҊH��p'��������a��������H��j��&��_r�=�������V�'Dl����^>��a�Eҡɩ�����pu��g�ekaݬ��χ���Y�����E��{���	X����<�����D�����F��@M��Ŗ���eJO7i/���������}���Pp��]����Rec�ڑ<TO֋�������Fi�r���Y��]y�LFI�\��
�QX�$k�|S˯�0�j�L�����d}`������כ�#T,՞�!�D � |v}�8���"������΢�NP(10�wU��Y�C�x�a|�/�ÁV�:z�6�� ;l�� ��گaƶ>�TR����O՗s��>��x��e_GRlra��m�����
�������71a� �$o�G�#�B��O�����N#�ic㥣(�]� )���U�;gQB΂=٪���V�)�� M�o$E
X��e��)�I�i�Ҽco�a�5���9;W��۷���O��Z�U@�H����q��2��$�i	مX�� ����R��2fz�ro�@�@�~�pގ�������S%n������52�45��G-(΅2��7M���R��-�f�C*'{�i44��Ő~:���c��-�NSU�����������/Ss�J4B�*%5��F�2�����5M|E���V���ܶ,�>�Xk���Q�pd3�`��9ʪ�������*U���N�כ
Uw4|ǰkF�z1�ƹ ��뢨��qC?�� g�vQ�8(B�f���4�M�)��l<�MS��V�	�w�`��%؆F�C�l�Z����F,�3��J��D�9�	�v���d��������1����d%��R��<B�`�O��l��S��l&�uڣ��������O{|T�@�����R4��j�~�7X�s?����K�)�h�����;���(�i�
5���5k�kZ���ԯG�X�;�Ͱ����沍ڻ([4#��7D6CT@�Z�1����T�K����}���w[`�ѹZ��"��^��{߱b�5h{�Z�^�ݏ�!(oh����q�m0v2������ې
0��m�%��Qf�(��`�XB�l�iG&��)��G��%�:��ίVlʦ�y���y��v���NY��@���v�Ȱ2�ZI��	����������ФK��C[)v�� UW$�|(�U�U{�s���49�h�"��zC�ޅ��x�?�y���+�迾T��i���}�ԍ�,�K˃�[ǽ�3��o������̻p����SuZ�K���\[Z[�h�%�\��TM)*"�TV{�M�|	k��S�<���t�������'O3�r��X�=#,��p�=�D�	����	}�i��*��,ݧOjS�b/�k��K.B*��ⴘ�"o�{�aQ�k%͎��P�X_=	޲L������U/�վ�u�Ph�m~1H�g�^������_��9�>��p{��:[���o�bBxZ�'��`,�!W'C!s��yq�\��I���R�������ıK�$����h�S.y��*Z_۲�L��ү�d9A��5Fb���Â�}��&�@^X�.t}r�t�U��"[.�8,���DkĞ�2���*Cw8�F���ڿ)1�uoU��-.��fi�d���)N�N��r�w=�9Q�bZ�C5&@h��/LȆ�b?��_���)�*�ψoy�y������̈��r�&�S����t��d��ܬ�kʼw!�t��T��M�V�e4U��k�G�`�\��ֳ����<Q���2WX�><�1�S`����Hw���8O�IKOO�3�$�3ΈW�~Ŭٳ�ui<�(IG��|��X�G�\$��XP���{t�|���H�y���>&��IQ�u�_���CLl�a��]��ꪋ���b`m����:cV�[���:�T�Gņ�r�`����Y�"��>�f��QX��+�=�P�R`\r 0�	�>f��{tWd\��!܁���7j�M��8�N��7���QBη 4Xۡ��Е�Kհ��G���Şm��4h9A�����P��I�v\j'7��`ӑ/�¿z(x��WȂ{%<û\SH���V�;UA�:$�?)�V���`,�7��m�
]"��P���~��4�~�:+�KQ2�s%���#Df�%�7G�65w�j+�QO&��F{*�2��_�PF�kG���2�+�Yfp~��1�k�'RR�#z9-ʔ��$ \B��W���k���C�J鹜%4'�'����e\���]@Z���^�\��a�� �uN,�$�r�F_��Y�va8}���v�n�J~(N{#`�z�` � �f�S�Ȓ֘��.ܹS|u���iē��CE7t���n~�4G�(�W����%_�,�w��+����D�X',W0��̗\�y���)l�0�UЊ-xP���XlxVHYEB    fa00     f50���� p8�(�O�*}��EP�K��J�$���(�)�n��T2ƺj�������\�r:�'[�L��ïq��\t�u{�T!pW�b캸�/H_�r?(�x�ԍwH�
č�)��۵!"K�O�#�8���$��`���6E6��R�6�x����¶Q�)�B�d�����j�ʿ�Y݇?���z�n�UĨ5�o�rgz�5bţn�4%	S�į����1�@�<�)�@�:�J]MW����`��Ȩk�긤��a���
�w��y�������F�3�N^����65�sY���6z�W1���-ho;i5s
.-�U����ڴv�?A�.k��͘�2Mã�l����a2�{�!�i���)��Me�&�G���L���.#l~�p}�c
	/���w��3<T�TW	��Pw�eO�&�洘G���A9}q���틬�%y�/��E�*�����W����b�i�}�o��	�ׂ��e�o	͕o��}�bS��SK���5��饤��ų7������(g��s-MMaD��\!��ɜF�.?��Ĵ�w��!�b��L	.�쮨h:_��u��i��!Bp��f�|�My�\�������LV��~�N�B��s�_�&þ۳vNJ��G 3�/Ϝ�Pɡ�g#L���9�כ[��(����a�ԙ~_#��#���c��E
iЗ���?,�u�U����3�$<�%F��Q�L��
U ����*��`r���ef��Ln#��CH��!Yp�-̟�!���|���
Y�|�>De1� ��>І��	�M�=�R�%rD�Q�����hb�OI�:o)��5 k�%s��a��ëL���z9�-H��<d�h��l%�6��Ň�P��H�
�efl�l��=˕ ���MBc]�lA�ó��:��ak���<x:�3������,��X�BQ���]�S(r
��,����c�{\G���f��4l��f��c�5������ߨr�t����C�lr�zmS����h2�4�Q�Ȫ�&.R'��ۗ�i�>�G��$CU}���WK�R\������o�/��뺍��D�v�pu���J��]5�����t�֒#���H��m���|�Y���X�u��{߽8���M��	Y�U�ť�n�+����`&$*�ؠx[����k�v�C�%(��ȥ��par�����7ׁ�5���o��8���� �2�[�Z�$V$g�]�*g�%;f��;����-�]i����X|pZq���{JxiõV��V����ZK㸜묆��S$�
�?Y��p��hhўZ�)R׫���L}�P�؝p���Q2�ޝ����NS�/u��
t�}*� ÍV�#S��w
_|��= }+˾<�u����A͛��A_0H�^�x��ݵd�[wK��y�'L|�V�ڠ�>%龸���XW&�Lb����ݨ�9`$IÞս�j�;�|��ߡ���B�AY��Z]�̟x`4��[��2��g�@�����AU�íh�|��d��a9ێHdo�=�� bnE�_�ћ	��n/#����	��w���;շ���2�ri+�@����_�rTV���^n�c����P-������(;J�7:]�&��O�0�(��������^s�Rܵ��������Př��sP��  �ڊ��Z��t��q�e�.[wt�m����[�]���!YC\�M�J�s{>W��J���25��Q�g�L^Nٍ�$7J���GNY��+�O�u�) G��3��?��7�.G;?N�`#2�yCm�du�w�.ɹr�����y��ZH'1�=Ѹ��(�&B��^���<���m����'�����O�r�������z}ʴw�Twږ���dV̯��/К)����d#�����`��(O�R*>�ab������y��61��[�]�ᚓ�(���Pӱ�D�[��a��s��!��	��|5�}�����).|] ���8���?q��W�)����4+�dQh�̯e���Z�o���g:��>���\����bՑ���HNf(m�m�_.�ʻ�d�u� ���;���oU&�5aK	��О�=R%0Vy���r�a�������~��A��H� �!V��-�:�odw�{7�����V��춈�(w
��:�Pn��t/u��Ez��R}K��^@�#D�2�C���Җ$��fῬ0+5P��N���N��̃�]��GS�|r#p�m�����<�rdw��F��öV4����d��#=/~I���#qV�=����o�:�q҃=�~m Q/��߳�=th���ykCb��'K�M�X��������m{�:��l�	�����+fo�&���'4�Z�ccT�;%�|+k'�a[o�-l��6j���wv&"�2��
X ��!"U׭ӛk�zY�ń��A+���$��	��AF`|+Q���XJ���3՝�H���j��#_DS��	�(?٨T-��nC)(�(�m�g�O���ٶM�Z�!1���W�PJ�7b���(�Z��*56�4Nw	6ir�ȣ.���x�$�Ҽ��r�U�Zj�?wN�U��0m�0�x��|��=�y�\��e䷪�V	L��k,��ɴ�?��<�x��&�+矺��-/Ŝ����cL�%R�a!���X 1K�c�{eT�s���S�E���GnDc_Z��j�DЉG�	?�H�&�Q�����)&Ba�.Q�'�[�$�85��v�)뎕�O5�C��E�[�?m�J%�P{�z]��5�u$��=W��⾱9��C��N���� �P&8̑oO��~&j�md=�@��DʅΧ�좩)��6���8n�:��$9]�X}l6w��3�<|���.���rC8�� ��j�}~n��Us@����o6fﴬ7�sקWm]�m�a�MR�~�g�K���0rAn��4��=<>�S�4W���b�`)�����&�.ru@jM����xM��ۣ�vd�	ySs,����K��t�'�G�S����~\��� FY�q�@V��a5xۆi��+��妛=�EU�o�Q%���*��� /�Xj(�Ἇ�訞U����D�܂ �ᚇ���ӕ/�l�Ś��ㆱiKp� ԑVƲ��=Evl�����qB��!�rs�l��/Z!3�h��}��5�X(��{q�+��Y�ӊ�>�-"��m�ݾhc2�Q~t�s� �S�[7��~��Q/,��]����Iʯ�L`pm��Б{|c��{W�q�
�V����
����hI�VM��f�bg�'�������OY��O	�߿^M�����>�%�}��8��h��6�*�gE�`c�?�Rך�F�j�W���P�	O*�>�d垲�����͵§V���қ��f����#�!�1���G��h�ɨ2Ѥ�|���#��R�(ʰc~ov��xU�C��(���a�fO�}�M�k��p�rq�pn'�⦩�8�������	)������=�V�T�B���23ˬ�?�f|�$��o�G�u-a-�"B5��+a�:Fw�H�Ʋ�3`�ֆ<�O�1\�XG�Q��S�Q�P�G˗^{9M�0rD���
��!�w����p��>i7ʷ��y��ؔU��?�U�N
Ձ�Ԟ��rG�ĕ=H�L]��#A�j���}ճ,��{_t�t�>��� D��Fd@|DG~ĵ}ש��wp��]k���2�oYG&��a���'�ZTUDBc��7�"�BI�I�z5�?;���W!�*�#��_�0�g������}�L�,q+�6̀B!OЄ{*-*�GN�R�6Z�م�.<\��FXat�� ��9Y�%����!�\6�q��Fm�¨{ >uX�[�������b������
�FXlxVHYEB    7273     560�t+m-s��P/�}�)I���>>tR��G�_{��prN����p.w'h*��d-�ĢIR�U ?��*&)��0x��D*���P�"�s��ƈ6��a��:�E^UgTwM3m�>������o2W������p�Kd_H�Yl�6���]b��4��|�B[��~���xćr���d�y�U�_��Ӻhm�����RXMH�adG��������c߽,�K��嘀���ȍ��n�ڹ�qB��|�^��� f���efvLaa׭�CM<Txb��C�� l]KZ|=�KӉ�tZ]�Ȁ#B!Ȁ�Nh��Ft�!�q��2��V�l97��(�q���qM����zH�,�"�&;:_D���84;ɏ�����eїĭ�{�=���8��j��*��/�h��ʕ���@��8A�P�Xee���(o���􇨁�kSk��{7�Z)B�	��G������Y����6��&�S�# 1,m���~����W�*�+�p�,_r�z��y���R��|˛6��Ӵ�s8o�U~Ӳ���(����zW������8�QT���/���9�̂�H�J�����-<	d��io��[���D.����P$����6]�}��ٚ#�*�v��f����۴JE���9Y_U�6��������´!��<��dT�8�q�\,��t�E�cQ4�>��[M���
�F�����|Ey�L���)4�Uy�
�c�:��G��&��7J9E����;��0�L6��^ͫ�s5���-qs�>r� �<E|�\R�G}����/��	)[�b���\>���*0����6����Faj��&@ܩ���Pԑ�Km<n�j����!�J���v���u�hr1B]�l==f�]]X����R�j7m��4�x�Obc�jGڲ��I�0��u�(Q�|��	�[)�����K���-O1�����-e�_�w-�D�]q�RNJ(!�j�T3F
��	��<��y�y8�&|���M�xQ,��U\6�����o�����Xs5#U;�Y��)�^����Tc��_Y�6���	���&-����h(J������^�����CFǍ�^�5V�Ӈ��A�*�a. V:6��Fw� vY
������^LL����4X��Q� ��"wZ����t}Yb�8�x��<[�:zT��bE���-cq*����X�\�� B|�MR�i8)A�/�X��0&Z��&dY9J����2X�$��
�#&����2[f6���$�����sY� 7xawl>�S��� ��f��s��3�^;ɚ6�=n|	�� =��	�� �0�c�7�&6?���Λ��������<Jt�A^ �G��;�]� q�6|�v