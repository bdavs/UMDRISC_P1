XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���fyu��8u�����=��d��ƎZ�d�z-�*H�oPe0$@�1��2H�~��^��e���y������$:���qm�����ތ��Z�I�U�Bw�m0��Q��{��Z=��Z�s�| 7�xAw\�D<&����e-K^o�W�����F�����7�;��@�X���p��dp/�67/��a�������U`{X�)�^uxG��S��A�N0	�**��JZ �H�a��[�L*�}&�E�@�I����I{'֒>�\I���e��/��eëk/�'v����篪YP�b5�r��<B�(��u�t�y�dY2��]�7rn�e~�4#��'�\�d�L;8g9���}�=ZU��Һ����H��ؕ@�9qT7m���~�uƔ���L�ң�X[s׺\�y>����^���ɥk����E�_�[r2�I���-���ӆf6C��x0�V;G��J�a��FD���hBx���R��9�z��5��uߍ{��
?r'�L�""+�B{.l���cz�d�t"Ia���[p�\�����!�@�K����&E����i}����ZV�?uix���t���*�X���Z㹄��Ox`@J��h���)�KF�1��mɲ��$Ύ��V�p��X�З���U��3�%�,-Q\e�ó�����o&�^!eҐ�Q����0NIG���9�6b�]�*Z�(���-�f]��/�n����^����ԍ��#�06eq2m^$L��/����t;�tz�GUXlxVHYEB    1427     840u���K�_	%��rr�L�����o����#����&��[��B�� =����uVOS����`T�!��։�G];"�yʔl�_�������|�H�/�)��۹�N�옍-=�J�%ł�"疠�}�?ͧ�,T�J��}O�]�3��ܿX'd&�j"�ǻ$P��S��y�5-�c�L�FM)�A[���':4S?�k	[�y�f/;"aZ%��4�ov�9�6����a���y�p����� ��	�>�'�@�TAq��X��¸gO�Y�jm1���\'��6-�3y�ż^�%:�?@���Md���Pe�r�n&�Q� �~gz�L��cB���������XڏCS�zH�|2:�2(�t���׷��`�-�ʷ��Q�[jk���%�z�O��i�����h��ecf��	S�8.!#��1��_�8�?�S�e�M��-j����;	�����1w�}	DT0�Ga��ȒM���N;s�&��Iܛ8K*�^�)��H��e�x3����'�;�3(Y4���w�5��d�g�� �����~J&�_l� �y�[]�m���؋������jH%�ClT�lU]�׃*4�q-������ �(����O���E��ؘNIu��-Մ��'u��m;aj������%�!)V�ˁ����(���O���.�O��`�!�SXA!���KϵO����[9����P�T <�'Q��oy>Ys��AQ��!7*פ[Q�����U&8�^�v<j�Z\�y��l��7��(�x�VU����1�v�7��ќ�ƺVv�9W%�
A�=�Y������K��li�$�SN�@�ý}�1��r��▙;���	^�$}��a/��ّ	A�(B;W��N1u�C^L��\�M����� 'WMq�p�M^���_��k
C���Tь�x�4H�a)xMV`<e��� ��&�W�Q�j
JRu`�#�2��r�I�289fHDH.hf�q�tw��q�^��4�eٯ�.�g}Ȣt�C�`w��w���JG���<o�d�e��Wn9l�(�Z�DH#�4�c�y��Ez���cc�H�خg5J��_�-��d^K��G�t\dO��A*=���!�����^�� 1���+B�mͷ«ß6ÒtQ\��1�e���a�>vc��)�q�Rd���[$�����h5�w��V�D�~IQ��J��xR��*�/`�������WUF'x� �6��~�i��׀"���,t�":�j�ʙ]Ե٘i��Z5���w�����n�%��K����o",��)��1bm���	��ߋ{��% �,9��v��$!hg�O�ce孝��A]�"O����E�? ����e�'do�K~�?��?�`_��g#�u��Q���n%�f̀	-��B�>CAV�=#F	/L��z��Fv�����^�L���-Dd�˾..�*ܝf><yLr�z,kڍ�1�~6������,���$��Le�	�F	�^�EA1�};�q�r�~�ͤ[[�si -mR5+3f��`r�#	�f�����̇�z�}�֚����OkR�Y�����Ǵ���E�q��w��t�y5	Į�(���Ӿ\�`;9^ԖZ/��3cD (�G�-�)���Z�G����W�D�Ȗ�䘴3�'Ӕ#T0���|��Ti,�J@�����d�/����g��
�}��bj��N��)�2�(�����;hS����E������9��+iv��=\Z^)n"'��.�+{@�˳w�ӂ��A�t��PJ�3�u��3)�E�&���	��>zɁ�)����ɢ�Ȉ���Ba!)�����%�����9�u�!Vo�W긌�nz{%cɀ�EE����,9Շ���{�H`�׹nN�c�ZU �'ugs0��~/���(7Q"^�!�&�2qO�� �`?�ݝo!u�A(�i5�[�9��T5���=���l�i��;8W�c3|pᠿb�V��i
��f��3��]=��x� Gb8E��8�R�RZ����iY�w�_ঠ.�"��[��c�yi���iz��8Y����4�XM@.]E��Pַ��{��FX!mc���h���=�