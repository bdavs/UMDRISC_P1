XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8�T��we/;r��H��l��jd�//�'x��U�Q�7,ƆL�Z�R/�Q���Nc��;��-�3X}��[j���y��~cQ&Y%�p7nҦ�+Q��/��=��(��P�c�Y���w߱g�%U
��u�V��c"�yh�\��XH:���1�>!`�8H~��r���48��{&����	��:dzbiFc ri[�-��b��x��ˋw��m��7��P�ǔ���f�'0A��bepZ����6��ro��Z�
Á�$����$�y���FyE>JS$?���Қ�ҟ^G�����Um]�r}�,^��sE\ޜ����Rf�8
ֳ�R�N���L��=�{�:���D|ո��=���T[���4x��G�X���LJW��A(�Ч,��C�'��G�ˑ��j:�d�PI��M��	!C3��&�%�
�y�0�{quM�����q�4e٤lTG��q�},�i��X0�tՁ��5=oV�^ mPȎ�p�p�3�m�w�S�A'�����ʡ��%���f��Q�05�����C�1F�����X���W�jt(��|�<���[6���Rf�6��ɠ��]���R'ْ�%�nd�A�v�1� ���T�y��x6��}���>�����1��C�ks���7��,^<3gC�$����1{1�6��h�r�������Ô!`�����P�Q9'��E?�������Ě��ni2X���n~��u�!h���)K�[�e-��^2 B�s���XlxVHYEB    fa00    2470+�wv]���+>H��f�N���� ���Bp�:]��_ላl��H�B�"��E��M�O94���Ȗ�GѰ��ʋ���麚�}Nw]`m�-(Ɔ�g�Ő��ו���:ׂQ�|���D7A+ ��w)�,�`�D����W�>*D��9�vQ��>�c�xh�)� 7�0�"�3wܹ"�h[�z����7��ʶU�@��#�?��|C�u:��W���棣����X�g)h���2[G�-m�V�2sqdT28�s9N溰f�5i�_��b����k��e�?�n8{Oox$m�Z��Eo\��݊ZGz-�;|��Z���>> s9*�9G�����h���B������v!�_���{��A0���9�E�����ۊp���ɞi�a�����{!	'7�/�� ��/�ia�3�%~p�����'���[ܬ�"�e��)�@^�x�N�T��k,�u+5Àu�@'#�@�5��,�/f:���U_ �+���pסv1_���U~��(����5��$�q88J\C��"�ۄcR�u��9͘�����/��Г�D�V�ZiPع�<F^p����<�Ί=�&�Lf{t�����\�r���Q�/|�e�t��tz$m�_�S���cW�W��=�iL ��}yY��Nw5w��y�])y �,2�:��)�E8pw�As3����p���B<�x��Q�����͠6mw-E��v�}t��-#��}�,�4�|�e�:Xl,�)�y��!���VB{�xx�y+T��i�s���?��w(�뙞o>�N�:�%�c�����D;��N8},�d� �:pc]����ܸr�R`6Q����I��/K�ע9j@�'/�=�f��k�]��J�e�+��f"(�C���Q>�W}E���Bg�dd*�D���"1��o����eM\��ww��P5G˵ be�\��<�N�nH�vu������a\�
���Z|S��Bek$Hy��R)�Piw]���y�n���Г~�����a����P2Yw�+[u���Q�U�ufT��C Nwv�!){�g?��+|�%�0�p��)/<� N�#Aq�c}��EAǸ���kz2#T1��2����e�SZ�*&���zbn='+��N�A�}ؽr�s�4�.ґ�(�H��Yq�qN���w��tP��&������ց�T��I�34�=.�wj��ױ¾+��u�ﱥr4LT)5�\���#��|�C�O�`c��K(��rP�v�LD(5D��W(��z۞�v��<&n���*��?��(o��=zn�?
az�:�2����t������ܣwݯY�Y����kǤH�������m��ǽ���1>��M_�+\j��Ex%淈�((,o�����
{p�n�	�ޣ0i��A�Ŷ�I��Q!gou��Op9X�!��^���_�[��*�$�Ń���� ��MUp�O��C���M�FeIq�O$[�����.�Jp�Td0��5g�y:��gpo#ƗQ�2Q���QK�/������nOob���o�.l��\����	��0_8�d a���!�qT]|]�O)b�b�N����d*9	RN�&��~�
�5Ϭ����^[����=��i�Ť�w�^؛^R�ؾ�ퟗ�]�}R��Ќ~BE;A��ڽ���,ڨ�؀��P0��n�s�>��� ��$Ibzmm�|h3�|�x�ˏ^�MFe�9�����%��b����|�㻂��,���(S,��]+/j�˜���r`~�f�1�N��z��|z{^�G���G��y�,��%z�����y~W��J�1 ��ִ��I#Ú��y�� �Q�ׂ�K��l���u�'��Q����;��M�����̔�Nj,��*�Ɛ��
�Wl�Q���1��q�cC�L� �b	^�����������R��U�M�!U7�{���<�X#@�?Je���W`|]���z����W_��Ld:�̩��K���=�!��I��jX_feO0=DF�7G5�6'Ǌv��ZP��~�t��Ȇ����S����U�JGE�8��hÁ�w�<$��� ��orG�i!�����ئ ���XdP��枣���ga���$����R<A� x�J�eW��B�~��P�4��:\���;o�6o�J�+��8�����`a�����3��ј���8�P�h"�b1�ŷ�]�����8Ng�?:s�˅)�F_�>UoQ�O�=�\��)��	�]l��1��
/6��i��=�L��1�^����0�$4ZI�R��n�yT9�N�9����ƴ��3����Cn�o� �Օ��&S�=�\ē �W 3��IW`��26�I����	��J�@})�F�c�f�x5O�5곽��j�4����Ϩ�w�)=��N�b�
�J��4V�tdX���g{,t��z�TudO�����]%12�T��b�����Į��<$j�O��8��sW�D����U[��1m$���e����nR����ԧ��i�����y�3{�K���7K[�ژ�]6���>xC�C���y�+fރ���Z��ٵ$Ka�j��{�`��&�+����
 ��ޮ@$��er�����ݣ뱦e���i���ip<��:���X����>�@2޺,lk?�w�b@hпb��dÊ�]���:�7���]P��r�$K�����ol�H\����sK��(4L��U���5J�
:����2�$dwl�V��^���/�Sf���9�G�h�t�8܊�-���y�z
̣�+�ͦ���q��1h�a�_��D��ma�K�ki$J��i�iTL����ex�:�� �ȷ5��
t�*�q�Z�������LҨ��ލ� �Y�ƤH�'c�1��bԅ�ߵ<�
�8Jw��v@�:n��ʟO�vȓ�z0�(b�-`���<���QS�h�g F!Ѷ�C��M���e�z��tj�
���f��B����`Sg��`��#0������K��غ���cp2 }��i�-B@�8�Y[Q8���D �BfF�C����T�'�)No)%��w(�}u��s�nS'�ɺr����i 'D��q���V���'#J���8�e6aL8eσ5L�HM������PUgG����2Jp_��Z�|�*;���)��M�w]	��R17x>�����Tu-��I��{(�҈d�y�e��+�b�5��>�E7 �S|)6�M��,@r�������<k��ۤ�=� �ß`��/��Hi��׋~���rb>To8��rmһp´qbs��NI�v�A#g�E�8ɋY8�ԷI�O��Oe5�Z�CWI�4���)I�ύK���J?6+Y۔e�C�mI��u)Ч30{�fD��Qu/Q�`(��P%�)*������	�j�9M�|BF<��Bz�T��.�����uS�ɫ��kg}f �=�K���I�����LƝp�F���'�UG��9��kUwn�y\<W�d�W�3ȧ���C��I� jT�X!1F"��|�dz��_�;�M$�yz�z4��a�h-6*]����HFѱ��f|b0s"�V�: uK����s�Q�_'2/c@i!�9-�,H�� �0F؍��N18���^�$\�m�?c���	TϷI�x`�a�E�2 ?� b����b��H {�59�b��@��HM��x�-�6?˩P<��1�__�~h��A�y�ר.nY1|ǿ��S��mF@[ Au嬀��pkl<�6������BS��(�VU��R�tkWJ=1='&�o H(4m6���9H�$�idi `+؜Dg�����}��%q]/�'���c�ܕ��9>M߀���ل��a��#�o�ɝ����~��Xf������Ƚ��3,��<�u��ǰQ�_?��?\�N�Io	�'GB���{M�Z���r�ҍC5�Nꅘ�2#M�4f2���4bq���KQx�G����3Û}�2���C��v�+|�vY������p�+ ��R<J'-jks�t{9(�>O��@�ӷd%L�:q.2�5WM�H|/�����>�����{�@�C��,d�S^��tM3$��w��r�,Lr��5n��vj�(��������2�O��mlx�ǽ�}T:��1�r��܂��:���]$J�T�n>Q�Xc޸�2��΃�w���{?�5�3xS
,�od���k���sx1�I�E�d%>�NѸ�3���p�;��=���u�0�]q�� H����Ew2x�d��ҧ��(�6l^&�� ��i6����c�_6���&c�X���{���I��M:)�Y���.��~�e�'��?^l%����	ĢEY�U�c*�7_�c����.����	̗�{�9��Q�7.M _ʽH��1��a����U	NF��	��RU�"�G�S�v���{�P<t,�7�WN�2`�k"(�Wc�6���[�ͭ�=WŁQz1릪���w��ѝ��a��XU� 9.��:�һ$�I�m�qnI`!:O�ׁ��'���F�uD����o;D��`��6�_$¹�j������ �O�����`8u�
\���x���Qw��"O�c�� �w�O��(�-ޫ�����*m�A�{�}h�r^�(��+���$�drL��8�+}�aQ՘�h�d�l�"'H:#�ڡ[*"�,���'ِ��^�;,UNV���gf��9��훁3�~��r�s/[~���Fu~ZFL"uF�Rz4`W�IH���~��N5�	�u8a���i�OHQ*I
.�dՠ��iFo]p��R���3�;^��DzJ�)>���B:%�1�Jݸ�|�E���k��w��M�Q]�T*��6:%����3�O�0�ܹ��Z�|�|�1�03��4B���Ry��+����_ ��}H7U�3N�g���՛�+��/��!y��ic��e�M0\1��h�r&:�1%��8���� ���ه�oQ
�Nh}���_���
C��tl8� �P�!����FhM����ۻr�D]!\b��'�x�<EF3�"�T�:^.�o,Sޅ���>'�Yʡ;ةێ�΅v�#���C)�`�-������Jx�s	J�P�k�$t"弱Q@f��X{aP�"�E��n�Z���b�?6*��|�U���'شRR�Qp�\��c���i���E���'5J�w�씑uyw��"#� �`�k*AfZm-��e���h��LɎ%��9�".E`s�(Ϧ�աc�á�^��yM�x�a)�n'�#�����U�C��N�B��*-�̄�2����vjrz~�����5"+�뾝��f#'>�x`�~\�*���ȹ#�#��[/~r��>����lb���H����w�QҾ\���5�R��1m�U|ZQ�߰~���/�#%eX�=�ƨ|�B�r�%i�z�T����x�#��������%$��������nk��m��|��b�$���o����ޓ/x�@O��o�YGg�G�ȡtg<r�W��S���m0D;1r�o�('ee'X>$W��Rb�iG�z�B9��I�_�7}��k6�����Bw��R�FC�ԳW?N�9y*�^/H�΁����u%��B��De��k+sQ��I�#r�֨�/��h����1��4����$�%|�]��8c6�-�Cfv�Lɝ#�;��E��+ ���xذt���U�A���B����$G�Z��TS�(BH ���5z�d��dw�_���Nq�������5{CNh�;zV���'����/į�U����4��U�����v������t��kj�i�ߞ
$���מ�:6�ߴHY�m�M��ݏ7P�w,�}����e�L/3�lv�Y{��p���{���%�x��᳇��>�!n�l&� ����V��"HǇ�9[�r��BWu�"Z�ʐ��$���Q���-�-��m1��������w�B�81��#����Q��)��Z�$����z��p�����y5[�Nm� ܞ�zc<;`��Q�3-���+�Z��<r���eꧯOJ�}��[�_�Ǡ�W�+�?VM�-3�dv��[G_�ʴn�Y�
���v�A H�K;�XI�p�+����}$m�P�1F�#����-g
��)�,�Tr����zl�R'֦��I��b|H4�#��ܰ��G����i�缶���x5���_��C��!;�'#:'�>�!�?������$ʬ��B�S�3�|{���E��ɓ���3m���0.r��t{`�Na����#z�M�zt"���-��C�
�?���8�u?C�n�N���iDg'd9���5�l���b �����P-U�λ5����]tS�5Sj_F�M�'���t�p��|�ai��~�9�O]ny��;M�f��~���:��8�H�~[=��J{��g�>T�ޭ�D}����P\ǠCs��i@��N�����<�?A�:w��B��q����ћ���|�Vn_�3ק=��0��ɍ�@�B �ۂ��'"�M�Z�鳅��?���I����t������Ai�|��yL�*&�,2�L�O�A��m8����>LBn[��l-?M7Y;&�D��mz{�}p���9a�p��Apj��0���ebYJ���0,��u�.�(��5Qy�Țm[{|���6��������ʅ3)�g=�Ë(��H��e��'��Q����0"WC_+{��e1��ns�C\��=��څ5��-�>X_���&�|�&��B�P�Ii���y}��1_N�q`�F�X�e���.���a���!R�OLB��DYǻ��)�.���?Y��ė��W���e"I���|��[�n��}M�0<����,��H|�^���H1y����f��&$ ��E�g��*�0��
�r��r�Z픬	X��`y�$Aa�҄$5z�X\$�{l�/*+���������m�WX���=��PR��y�		Yg�ޮc�����%�4(%~̐�}4��5"Ҏ2��M��Ջ�&��Fx�=\��ӨXt�=�C�mQ�\�wKqu3t�T��~�.�{`wٶM�.0+[��qcg�WwE�Q�8�}[���n�}C�s�/�R:�w1Y�Ȍ���m�"M��3e?g����]��/Z1R�Yf��W�q@�ᢏ��6u�.K|A����,v���t����)��ȶ��j�=�T�.���-�S��T�D���kک������M$��Dm����z;ҜK߫e���ѺV\.�?N"'C����U�p��0=
q^����3w��@ˤЧ���`̾F��y�q��͍h�[����$������W� ��`�u?m�����+���I�`����_�#���(��T�<�Ja�Y�ޥ�ڹ/Ҡ(��d��H%I!5J����K�ۙ�̚��ZG�d�}1wt)�A��]���̢hhc')�9���:ɉ��i��w��p_&! ;�іdD�;��Y}�}+�#C���|�,��i�K��j� ��+��ͺ�ގ�*~l�(���{� �
�ݒ<a�C�٢�,�S5`KŤ,�;%�HE�3u��Rm�n'���2wSv���.�()=׹\B:�dJ��{���K����ܞH�dm�=��T����û&�[83ckZ�R�<���Ϗͻ�w�z��.`n��3A���"^^Bҩi��USb楴�lf	u��yr;���{�c�k2�S��l�V���~�!&xۓ�&r8)b�~���$b����Q�ʙd��r6"�zh��A�9C�H���S��Ʃ�{	�G��r&eڊ���H]�$n���9J"���;$�E>i��>dS��O��:D$C��R0,��r���>��
��n��r�����k�Y(���`�QJ]r{������p� v���W=hr�0U�KQ�va�����К|�G4�&2��+�OUgGk��8��'�.!� �<7K
��:#.�Z*����t��	�U� ��u� +��b��^���4�L�D�Ld0��A'e���9R=�>���M����g*b�(�XY��ƿ�`� 'M��׉IA����kaW�E6,��a�o��]�j� 9s|AF�!_n
�6CHHqQq�,�Ả܅�/���!;���rs�bh��]��B�݌ !�p���tMc���B�se��]c�L:�Bvo�.�P��u�U��f���M��tR�F�k�����X��,��N$ۜ���7t���]MG�ٮ	��
���x?�!Ʊ�r�@ި|�<���a��7�o��"���� Wz(��k2@�x;�܆���u�vIx����V93?�m9[ՠ���E ��"�����q2G����Ѹ��h���5�k�_��3Q[�{Ю���,���K�V�k��-㪹8;$��� ����p�U��+���@�R�7�4�պ��)�E�'���$�n���;9���rU �G�݌Td�z��ތ���?M��?�\u1��_z�>���1�;�XJ�H��"æ�T�mats��6����J5�+��9��<(��RG���fΈ%�-V�d�(FJ�S��ah#��j#�I�%�t�0�lh[P��j�ƒwb.�iؠ(E�x�������bn�a��:����ɀ��y�[) �� ˮ����*+�0=<$���#�B�� &����s9k&���h󇫾�.�d�m*VM	!L����i��.�#G�����	�a�,�'�	�����?�tD�(~�}10�~���Qc�%(��$��6�stemJ����:5�Q�oyxC��:y�;�蛦^�GW����"��M]��������QX5�݇S����#F������_$�N�d1`��G4������G	 ��(N{�Ӌ�TH`z��O�כ(����˘p�1�W~$���_ZN��Zv���>�6s�[|��sv���ya�щ���O#d�F�(�yBY,n���q.搅�}��B*�/�%��[N)`Pjy���dX���T��"�{���&�צ���g���a�D��N��\��*4��)cP�"6���gK�xQ"���{Vrk�Z��N���WZ~�?�*��B����&�� ���r��"� ���E`�s2ٰz)���G�h����\�A>���{��Is�N��$C�*�0YQ{翔�D�G{��9�ƨ4�7��iUȊt�	Kt�D'�89�_ԁ��������-�`RP�n��c��XlxVHYEB    fa00    1b30����)��	/ŀ5�n���n��˵�W@2vZ#u�kWG���wP��tē�6G�
b�:j��i��Ș�7˥�ִ���PҠD,��!k��R/�c�[�RQ�vP��0����4�a8��@����u�>�C<'`Q��Řa��n�-�.Ǫ��}/׬G�H��\~/���PY$�BMrcҽ����E�m�ţ�)�}LDb������od��>-����F�|u8Y��b"�/K; ���xU�M�K�����a�XE.�V4���o$�������;ƣ����������f��������C?�b�k�>5��e��@os!v�����=T�t��N������ �0�:V `�"�����NX>��HόJ�H�*DD�	`��ex`wQ���w �boZ�S�=����K�fE�����$��������߱Ʃ$��a-Z��#���u���J�7�f�'E�;��d�:t-�c�W��A��itN�Rܧ�C:�V�=��9���Ψ�Јe��&��� 8�0�����ȃ�(ƶ����"��8��>���ʾ*=�5�5�I�8�[�f��zaQ�1C�E]љgT� �ν�Ec�(�W��9���<��,b�TӼ�iU�P���V����2L�`�,���b�Ŵ�]��4��������- 9c��}��^�=�q��/k'��Yx�\���l�[���s�<7��ʚQ���i������P�Ꞑ�"�K��2��#z�dx�E(%���i��y�K*?�?3$Q{;�A��2��,*-��|��)E*H5����ȈUW�LȚ�Os�9���t<!&�a ��ݓ��Iţ  =�Sd �p�(W����{bБmi�*��%�K�gB�0��g�J�a��CaU���-����ItaFZi��	c�[�p>U���9g��!C�(|Hz�n�Nv��ʏyN.�_�Mξ��{��/��k`CdE:�.耫 u��Y�9I����t��ƶp-!�VaA�=�_��u���sdK�:�>��u�\&�� ����T��70�6G<
~�>H)L�H�i�����M��%��_UΒ��)4K�Y��9�,#��:"�.��p�'�zQ+�\v��:�HLt�c�����+ n@3L*�r�$^\����X6�'-��_2n�a� �%�h���v3��P+)���:i� �V9�ú��>]s�e�̈́Fl6��4�b d�`����KLN�D��Bdz�����Dj�j�;��?+f�ϯ��n�B�ߕj�N�){�>��D�9�kJ���ڜ����LV�λuYƦFH��PH���/������`���6>jqf��S�ZO�(�B'VL�A��ߠ�4�A]h�R�4 Y���(�r�d^��Fq���*�I��~�׷K`��FH�-�������/%��͋X����cA<UrC������q#l�j�%`��]�H��|�y��va-��Uq7ֈ+ט4-��Ti�c�r˝)kWNT���Ƣl�:�@�nz�Y%����Q�''*�~ALߩ&��iU�K?����Ag<F�kcn��e���0w5^+6ѿd��?�c�0C��)���_�h�����o�R�ƕ�C�1���l���)��1�s�e�C H������7͵s���;���v��7��G��r����0���J)Њ�;f)�4X����l(K��6|�����Y����Aq� �hjp�,~!b�)"1�'v�"u���0�)R��`��m m��n	x��yD�b�sG�.W'�`��<��ӧ��h��x�z�n5	��0���7��̣n6�7A�[�<n� �X��V��R>������8�l=�斎���i��<��ldkJ�?�35���~��gDJ-�$)�<���F0-��rr����YJ��n�+STCfU;�N��pp��Z�1FP�n�}#�P0o�b/�Qї��x<�C��ET�%���L�kt�#��yϦ� Iy�z8�8�L�����y�U}���2���J�2��N���,F9F-��=�a�7�Y@0��S���6 q�+*��$�~�P3�u��|�[�}@n�aK�(;�pZ;}H�ű��u?����������7p�wa��`����W�;|�σY���U0�16wI����/�!�*��g�b��]T1��GK,��Ӯ���?r�#�Zp=� `��8�RC��cJ�5��\����g��v~�g,��i?����c�������|0�zx����0\iUWa���frS�_��qTS;����� 5V��A����3�X*�O0W�r��stC�}R�*Շ���;=2��I	��D�����q��w�M�SÖoM�2�"�5+�/��M�
���p�Q���YO�A1����/�=Q>�&�xg"[׎�׻k�w�2��/5�
jc:R��������2��v��Ή������vG3F��[�I�p9�R�[�E�v	��(�9Yk���m�lB���k�R��G�+ag��K������9a���޺LL2Kc�D*i�����'�\����uC�Y�Vr,5 M8��׾��D�t�E�W��E�	Ov,R���@�W�!W,�@��
�Mو���}�6.`S�����u��� g@R40�c�yl�g�[{>��/�~
+��4A�5gt6�Ct���L;�m�����h͛5|�U&�E�qӄ�����yV'.j����0�,֚;�4ʌӚYG�^�er3���i��vc��E�譃UC��k=�j,*�b^�~~�w�D��ޯ#�������O
�
�D�,��X`f��`!�8��Ӭ"�q����e�$n\�"�\�!�~�q��YG�X�."�-���b����o�d�X��F D�t���83�@n�oj�6���M��K�v�2^ސss-�74�*[W1�*�#P�j/������v����*Ã$K�+}	J"�Ҭ�h���������w<�z9�z#"��Q��>DQN����E��r��&��Wȇ��ŎQvg<D��)m� _�H�2��1��g�^�UM����	p�E}�r
��=Ƙ��=Bu�c�.�����?����T|�B�[*��z�W�b�ҷe���~�e�����3���=osb�3pQ�����C�s;b�+OU@#p�^���T_]]�(v��,�jxJB�̄����>��RDE+�+S�Y�$���;�,�� �lm'P�r]�&��^��៼�����'SJ�.N%Y|�Vj���u�=Z�\����'��֪ɨ�"K�=ZC}qK�5�W%~�T�F?of�5ik���z���e%'~�u�eF//���;�NI� �N
�l�3���7�n-�D�h���������a�Lo����-|���g����p�͔ȅ�
����+k��GGFQ	������5C��B���Z���P\-d^\�7cJ������Ժe^�6˯>āD�@�&�?�Z����+�\$�^��>�7�d4T�˭ D�&M��"�����t�,%���]��������$hg|G����5O�4݆���d��%�yk�Cf�;�3E�9����Wus��i�#���3HC�jV�F�p�#,V��������sopX��t�]Nh�8c�9_��~xc��.���y�aK����WZt3Ä�U*=��TC>l��D�4o�C���=Ȼ1��g�k�^Z4{X�,)Prb�ތ�+�K);�*��+V��T�߾d��L�$IL�*�e��@���3����������>����l׷��6G8�#[P��@�C�c_L�z���a�r/7���4��ɪ���QQBk�ݎ	qx��zvH)���r��V�Iv�-�����{��%�:�`�q~�ψ#M��eu�3bDToG`tVB"2�.��Y��?����j��D��2�����L�5L�4�; �@�B��?��k�EvV0��O�cX��Uz���':�{Q�AƔ �%n���� 3�+�j�Ƥ��(0&�����<���"�RLr����=0q�>{�����y2X����AQ��<���,�����}���	"��]/��2#俜w#2g��w��p�N��a���-�T�Z��M�5E���o�,ڛ���6&,7�����0Q�t��߸Z�`~f��/�I��5z3���Jm��#����(����:
�d�*���Y����//��̶�ye��Ȟ�M�����~�>�����J�S��ad�&�	;�����s��A�������p8�a��w3�n�nik\�3��>>t7D�f��M�uL8�&����ܯ/��V�_Nm�?����P�D�]o�Kd"E��ѽ�)�#ﻞ��C}j'�����) H��i��Ȣ�bܟ�ۀ_�<��҇!���V�y�m>�R����i{]R�n(�=T�C0l���^���~n����������[8�	\�C���À����\���(��ɔ�e{�c8�S�K�~��x��RoI��ek�i:�������F�K�D��Ƚ��{i��DV�t�jv�r���_�Ϩ��j*S?SW���H%A��������F\�J������L?h���AC��a����\��*������v����]2q�`j�����d]�_�A�X;<8	NX6�ux$7�&��o"]�2"/��@#�v�]W����o�P��%��c
'@/ *z
�u�CkA(�l�e8Z��v��E|5��R��YfB�-/yf��t�VY̒�*�s
��8#����j�������>�(�uB�-����tv%*.�S
aͽ�3��vqG�<c�'��Y�-���[9�oO{�=�W?�#�x�3�+-��k��̿V��Nx�84V�������X�{�#�B����'m�b��٢��;��c�=��V/������e�E-�q+���]�@%4Z5$��݃��ٳc�R�4�����>5�|:;Nw݄�u��QG|�yf���)��8''�uḍ�ԫO(��Tz��2fd>����V�ʪ!�^���נ}�$`)'��#��&��M]o6V�Jb�~���vO�����D�B���m�|\⓺��H�.=S½�[���ʱ?��tE�ۘ�x�2��Wœ/ �R�]N 3U6W�+��7hg�tM����Ѝ DՆv�t���A%�cYi
r���uw�rP�JU���HRE���MJ��D�9��BE���w~xN�^W'"G�
�����M
j�Y�%��kX�@M߱D��҃�?���H�\1w�߆���*_k~oԺѶ�]���h����!�F�3�a:J������ü�vuZhB��iH㊼0vG������2�es5���ˤk����	���^VOmA�e)H�[Bʹ����r����H�cIX%H'9�+^C���{��Lx�_�~7Q��&lj-�9�8��bĲt�ͣ���W=F^���,B���,pq����]�NW��=���6K�r:7�2�e(WՏ���鄧�"��]���)o�Zv��s2Y���$_��������������f�t1Gǈ�X\*�p�)5������?ə)��0,�o�u��,Q�6�m�(�ǂ%Ļ:%Ⱋ����6"�4�#�H���}�1!,�էd�/���w�EWͥ/�T��{ �������త'R�.?��U �[A�&&�&���M
�q/�}8�B&�z+V�?[ӄ����f4��}=����85@�%N���I���[Ia����c ��e�n�_�P�E���lp%�����zZ �p�7t�S������X�� �S�YC͋΢:{L��W��:�Jm��}Y��7==�F�
�z��Q�W�\�x���FlO��FC���@��_Z�l�݉-�բH��J�|: }�F\.0��<�C��j�7y�X��aph��5?����F ��\L��^́Fvp���m3O�ķ��.�)���JTӏ�=�IMe3]~HA�ޟlDŰ��K~�M�Gb8l����R-.ߗ�E�WC�}�UU���'�W���d��w8y=��hw	�tb�P8�)o�wx+�ΗJ5�)��X>B��H�Q�:r"츷�.�~T���#}W�b���`�IF��Zl�������]s��e�g xx�%'D�Ӂ��]�����f*�Y�%�R��	N�sl��IT(�F���s.l�,��ڭ�`4ܢ�� ��-f@�~���K�
���9�'��+�NP�GU`ü��!b����r�ӂz&�>���v�z�c%FD�ZBX��K�vV�UD:��S`���R���~�Jp�h�e!;?��;¼�ib��=^�ぜ���(��,t	]��da���L�͟�����C"����K�1BSX�9�q����3C ��v�[&�ȋ����S�0Y�Խx�����R޺Z���V�~S̥�~q�����ǐlh+���"�,�\No��%K��t���f[	W�N3Z��aP'�ވΞ�Փo� ���;/L�-�l��� ^�L�i�Ps���.�sq�|�ꔂ�K� �	7༾��P@���@�P��A�K�T�JjF#�M�L����q˪�ҎLCCg�a�<ͥI�+����$��qâ�����!6j��Xd4����qtA���
p-��y�,l�ʴhO
�W�h�ӊ'����
8��u!�F��������a�<�6���H���Ǿ�[���3����󀯚G.��;�>�썔9��a�k��cǊ��T��0T0� ��6�;��^��X���P��}�>>��8��]4��4��@L�����εwd���ȜW��|*�2K=�'H�<�,}+g�7���	�tb�T+���8m�XlxVHYEB    fa00    1950G��Mښ?"@�)�j���^ɗ�w�����rS.���3}S;�Tv��H� ���H5�$'>1���k��8�C�4L���5n5�D��Cg�Ƀf��R!�AQ*˫�x����"Ƌ���4��5���(r�@�zQs:Y
�B6X���k�n<|9S��?�0�_�l?���;�T�㔽~a�+Òխ��\�0���)�:G`+Z�\;�����_h��FF�)p ���ϊ��%��Ms����'#=�7��|Ғ��* ~����O0�'S����!Ʃ.�aI�*b��
��9DnDv���s�;�����{���I�1�<�A�D�`]����2��1O��X>u��	��V�s���f�\�~ӿm�fV��)�I*!�3��[�����vA�K\䬔�?����C��^���.r��c8��%������S[^��x��7"So���b�Q{�̬3ʏ�����m��Xd��d埃�p ���j����Kf�1r�?/}r�Y�*'��V�������n���LYU ~Z��h[����� �zbu���I�{�m��ܢ��>�����2����PgF��W��-M5�"�;��K������Ru1#=F{Y��F��Dz���B"�$�C�!wF���u91?�Nא ��>��,�yd�S�;�9ǹa+�А�f���㮭�ϖ�bd��fJ�m��s��r�Y?������dzt�S�Z���-��Gn���U��3�´h��ՙ�/92@�\�	�??���b��G�B�����FCKW�FIXt�$Icz-�Ǽ��;�ݦ�%�.�o�~����i�4U&�juo���L��B`�D#������>X"�Z���M�k�÷%�]>��6y��T�Rߠ�q�B�7�x�t�4=�}g�e"�pc�N �o~B��\�Upj�v�a�9@.� �|��?Z��Q�}��k�t��LI�W��;�:�W�^>%�s�}b����*���	j�7<��1�!j�З&�-�
ï����k;Hkn	tX�.U�<�	t��a`y�l�g�|HP�6i��ϋ�8���x�@�����4.��E��4�`�:^�_ǎ�K��IR��`Bz��p��]~�l�d|G �	����o���E�>R�zd�F�V9ֵ0�_gI;z���70C��mʪ�yz5]Ä��qI!���E녝vp]'���OΛ\1`�
 ?�"����d��\��x�;�	�˲?�|��D`0:��fD��.=�|��8m����!��fzI�H܊�7���@-23�^E����z�� �������p�x� X���7�0$�� ����K/L��^���~y�w�p4����2�_���)ݗXS��!��d�%�Xt4���Vϩ���ѯ��I!q�B߄w�ʏR��:�b���`�D����Y��Ѿ8&e��	|8�70s�r��U�-���g��oO�� �e��p>�FTs���9k	0�P��0VQ�"9%0�>��X�4Ld�jm�KqͰ~K��D����$G�����t����n��;�L!-U�"��c����$S���ď;[+C߾w�&(8.Q�IȈ����mj1���;�6�EQ��Lw]
+ګ�#taP#�pcc�K��:űϩ.>]�#������=N�vf����cbo���Z�w��W7Mx�H�j��j.,)X�"�^/���W�i���ؠw6ZHa�� 0�P(Ӫ���ז0Ne�i��?�I���'�a��k�\����խ<�y�ӡ���V�z�A}-�O�U���5��V�cS�����ii�B���I�Y��p�%��K#wԪJD�Ƙ3���4@)a�F{�u8��A�r,�۷Û���z[J�m5����{)G�+�ۇ�ox,��yѣW@��-�X-������3C>j���z�."��+�r4��P�N�D�9�����ħ>2�����	���֜��{]�2�b�_^��Ƒ���#�YL%�zd�����~q��K���#�u�@B���[�3�<��onJ��E�qm׌�p��޵Ga%��|��(�K9�ͩ�5��]�'xM�T��"���W�<����
*tai;�Ndأ��D�X�v�����Gr!��w����[g�_�� }0m*�D%��s�;4�`B��dZ���'j+�r����'"t�k	�N �'�~2�Іzqkrk�E�mD'r�
s1�0�d�~b�̕��;�i	��N	�p2)��h7)<2��g�+���(�)�N�h�^u�y+�Q�UT<�<���e�����,����%�Ow�h�Ґ9��e��l�sr� ���_���/�,A?�/i2�ң���N�����*UC������h�2�J��[Dz���b�av���w�4�l':,����[�||NEH.��i_���|IA��2�����F�s�D!K0���ieD�l>ſ3� f[g���[�E��T���[bMnY�Y���~$�&r�ɿ|�p�����ٺ[�*�'�9�%��*Y���=�<��	ψ�nj�-���bOb������;�R�$"XQ��ճ֑Xȿ�EZ�eCN+U->чǝ�I�b�[�UC�|��A��h)��=o!���
���*U��5K;qa�5-���������S��h���<.`�I�[A�"q.�˒XHZj�(⦋5WM��J�X� �+�>Hm���X�|��F%[�X��V_��GԞR4�@�dµ tӓ�Z|�0��G�ya<2���!��,ĭ�ˡa6��R"&9����:�t=筦�z?ث��8_�yR\Kߙ孴���2	�bɤ�V,^	���3�Yx>�d�r���A}�]e��^�D	Z�B�����G=��q�s������i��z��$�/q_�5v���p�Con��>R�������<?>�����3�l���̟m4E8���2������5��A80�%v�(�Nq���2�Y�q�g�!%��-J})|����s�b�\Cn��xݽ�IZݘ"�� H�S-N,�<\-b����E�,\Y.<&��R���7L��-1ʵ��I,�j�,�� uǦ��!7��AI�� ٦�3�lRxL���^�ߙ�}=��Ҹ�������ʮY��U�����\xM�������C)�RA����U0�[4Gֶ���% d%pO���6g<F>0T��+W���c���K���i ��7B����x�_Q\�����NMO�#}���C�H�|�8��~�������^L�;��,he��z�s�2(�X	ZL7��	VT|�v�a���2:B�u���86C^ n��w7ٓ�.�$����k�vx�eb�E#L�SVu8KY��O���^�vp�k�l����� �8(��x�!��y�g;_8�{r��pգ̐�o}��
8�P��˚QS(p�bJ.d�/�������5sw�>�)l���6���Tp�1����u���Vȥ������:��_�o�^��=4���������>X��-uF��-'��1���}�۞�>]�d�k`�4\g��9/9�5�J�B4��M�/�U�,c���Xo�"Whl��n���V�������f�ť���� r��
oM珓.����`�"Gz98#�SnYkF�oa1��VM����cM�$h�u�6ݓ>}K	���}Yo#�TKKV�g>�y�f��n�4Pô����Y��z��}MT�M]lT��x- y�wʫ�>�t��N�m�	�{���t'p�l�1�Z�d9{�.m�輣��^�>�fH�ބ�C�uv�+��Gc�ʝ��;~=Q�笛�QJ
�ٓcܓ/�$fu��
�|�P `+���RZ�VD^x�J�J4�.��%}�T⭵�wf5B��XjV���Ի��)�4;V5�eG�_c�Q�ˇ:�,ّT�҂ �����[v� 3KxgY��k��n>P"��h��D/M�eE�{��,oDrXxDѦk��^El�Tش��)��.ro��YÍ�̍�g'd�+��kXl>�c��-���MA����������G�O��x���7��q\���x��tpEs�!#�I���ow�e�#s�LI�\�g�ݛ:����8Urr�������j����D��{-�kPʜeG��T�@h|�6
��@�ZRW^�>�t�8��_����H����̟�5&ջcu��3��D�$J��;�ǔj��v�h����?"���]�U���%rCC�\S��!�
�ef�G�FA�h2�?!���^2��(aL�S.����$JP��.�w|g�
j�W�X���� ұdK}ޗ�C�ir ��I֒C�iW��䓑L�S�7C�s�RZ�ɡ�h!I4%�A��-��8������jۑ�����:*�ȿ��
�vs��=�K��T\.�G�gU��`�@5ش�w,F��i7�厨���C=i���\ȸ�8>/�R�������+�����28+8Y�������F�@=��9�'����8�y������ ���9(�l��s��4��P��n�U>O�ԋt�D��ôjx/�PP��j��Ԣ�=�e>QB϶����7-ݜ��.��<�)���d�SpX�ӻ�a!��<=�lP0��S�<jrD_�Ж��5-"�>R�n�l��R��/t׫Y�e�b�,�aK-a����<A�u%*��/B�U�=2�����+��n^� U�G�T�ݻHO�e�lT�~�*}fq��dˋ�`o��t�j���Q3�G+��6i�1tO���T�.�DbY��1�!׋Fī�,|4	���M�\�q5@_�x�)��V���p�L#�p-�Q�$J��`���Q�Aʙd)
����H��d�8��VXT�~fIz��I@�����=��i��Պ;#u�k�ߩ�ќ�1���Siѓ�!�u�Pe���騳�����E^2u�p�۳"��Z��h��65����K��QC�wbW��p���'�!�m?2|��u鿢@<��/��o�s��xT%Z�!�V��;�\�۝�I1iW%��Y�RZ���؆D�GF!�<��]���4s�o�q�p�߭��6_��
�ڻi����Q"E�	���ƍ����P3��j0���x�8����֩��3c���(�dꐬ\J�h��$�*u3�,(ߡX�E���
.��`�.&$,2���H��sr��e~��`(��iÙP�MbCa!G
���WG����`3��!U��U9��}�G�?|��DY=D���P������@��Yx�P߫����=<ϔ��[*=`�bW�{�R��!;������D3�7
�
�R��Uר��ߝ��]0�:���P�t���+#(�_�ǭt��8SL*��1�j����RuO�DQrA�\ོ{��(d���YG$W����������8����/r��j�pFA�Q\o|�����5�6,=��x{`�D�?�o7��j��$�`�a��W�@h�?w�W��VWF�D�������>"� �	�����L��,-Rs3j�+�8��K6'M������e� ��bI��3f����Q��5U�K����ol��������yx�*���>ü�N
ڮ�x
�� )���e�r	�D�h��j%�[p��A�P��B��U�]���������4D�Ţ�f�/4�3�B�m?o97��a�3�w�H�)8��q�)����+�1���s�A�}L�fV��ݘ�����Sx��!,�&�	K�|͸�1���z� x�b9>�U�$�L�UP�'�Hl�a�����ihrc�sQ��ͪ6c6\��N��5[�;Lb8e�l���;.F��w�����gU�bc�u{J�h�`K�ś�K-��2�`����W<Τ��Ԩ��b?�I#�a��j�>��۵�
 ��#܀�����M��������6P�ݔb♧��OBʰȷG+�4�J��-h��>���q���X���p� z��6���p*���+g�����I8�	ƋV�����B��TG�K-�KZP&{��/i#�L�;{m����]�(�~�&)�0�Q���x�,U
f��9�kRU�=d%!�����Ǵ)�`&Ջc;\�LR�
�cZ����	T=_S��Ϊ�l_}z��d8|�U��q�y�2r'��xEk/j/Cv7� ��a{b����?��K��;g��p|��4;Qu�ּ�q�}z֗1�[po@(7�h�k��K���PvF������(6E�ϯ�D�� 1:�� �\7<�>��#�׽Q@|')''�dA	������_&�K�n�ll(����:�����{�I��Z�k�X J��cͿ�I�>�@�96h7Ծ��"�2B7D��$�c��.���O�2h��jcCA׊?d���?�� �=*z���)�d���I~�XlxVHYEB    4f27     d40����|�հk�%%y�~tG�1����сm�|��t�����rQ��p#�.�`Ir���l0�.AUO['��B`2#%�\=$�M
e�}�ҟC��G�����_$§����v���J����<Q�x���P:� �|�n������X{J���Ϡ�c��F��k�.	R��Ct�i����v7�C�t�|�����l�k9�o���96pt��FG����3�!:��C{�Z��9�e/9�!{+�s��$���${Ğ^�`���;�N�Y�4W;�9E��m$��*��9�R"������z[_S���Xt������|$@�����|n����u 톹}�g+��+b|�����c��Q���V�U����Х~W� ��F�ن+��6 �e{��2L���w-�#�e�ꂂ���bG��:�Y&�(B����3{��V�88���	T���OL��ekZ�R��c��P�(UB	��(�������-����]8+ʝQc�
�O���3�^��V,�j��#�	��K��p'ޤ$���v�+}]9���?ф�՛.����M���5�|q�����^�?C1a�L���T�;��־1�M"#�ڤ��K_y�� u�A��c�r�5��/C���U.�q�?�Yr7*u��1;d�tzi�$V�������k�JC�OKH"E+>�C� ��`���nu�&uN'r�DRC���5�F7�s�u��\ɯ}1�b����N��Ed��p>Ûʘ�=��*}�_��a~؀�A��oq�n�K��)1/G�x��\��[>R�l�٭���
��]Am�z�ֹ�ϟS�/WQ,����'֊���.Ū�:���x�hP_�Co|@�~���H�2)������d7����-���n�ֻ_�Y���puD�,�{�2�W�+8_�.4�`�&r߿S 廕A����m�wD�����@�F2����dlʰ�,oM���B�qڴ�x�_��AH$n�-�,�g��T�d�'dW?�"+�H��g
i�./�� *� �������%����J#���_�4�:�$��>�N�7�W�N���9��/����iY�9$5(E	���b:��{�3�,5IVK���/3i��V�霑ZF%�x�Hc��k�(%�~ބ܈ۮ
�p�.��0�C=��od��f�D0)J��}Gϊ?���E�"p�v^)%ifv8Py��� ������i+��6��jaln���x��Q����ޤ��W��
f�t��u�7\�Nd��M�*%T�Y���>�	A�M��.����=��M�B���ȐC�R��v�����6�)��>���)��oV5��sha��p��xwB��q+z6��E��[ʲ��7��D���k�+�tf�P�I�V�.,��ūu�v؇���Cڸ�o��>ފ&ܛ�D�9����QN>�*/�fʕ��&��]��W	��i�و&q��)�&ͤ������oT�@���*gW%��pnw�b��rb4�@L�2v3>"E�[�F.7�p�;���0��&G������5�L�oU��_��v�U\[�Ok�RZ`���H*�{F���G��ΉGh�ZU^�I/����ڬ�4)�h�
Ix#��<a/�T2&�Ylp�� �� -,r�AS��D�M��d�jЌ6�OrZ��4)'��x�>�<o�8b�����U��E���U,}5U����vB��� �㊵�*��X	�Oτ�w��1��$*�G6���A��\���v��#aȬ֡��*kˏo��Ɵ�F�Z�Am�%�	x������k��ns�w��X�6O��^އ�qo=
�rKIG�d��	���J�Y�gO�-2=Z����X��i��ۨ��>s�����U��s�%��:�=c�nc[@�*+��9ZQ��a[��R��W�[ɞ����Kt�-����B]9�h����45���Η��X��S�[�0f2�%�rm��)%�}.j��=Mq���͗��5y\58R�B�&��ۈ��÷��/�/����2�R�c)��.�`d�|��ș��gs��(� ���`�F�.�w�Cl��h|³�*�'�xL���X,Dr�����:;0�y\��}u�UJ
�,��;GE~�ݣ�U#A��X���D%��"o��b)�B�t�*6��N@�� �Z�y�7�/��)}�m�<�#i�{�:\�O��'T�sb�v�R���嫪k�������&s��+�u�ϩs�MO���Tߓ�?��� �ҍC��^��ְ�Re��2˚���x���@0�Ϫm �%yT��:SL^���U��'�4����H�rZ���܆�i��5���֩F�qvgC��uǬP��K�Tb�wQ���U�k=���a���Ӡ��\�����	�5�tY[]��$=�9n�w}\0��t5�#"���y����?�v{��	��s칍S
Ɔnv���ńEs�?����-^��cf$��/I{�3�g��ĉ=^�.vp�~����Q�u(��i�扲C��3�l�/����6�9[���)��}=��� nV�a�4����>�u�*���T~6�g��yy�}=-_����*����&�eE!\r AH�tQ���t��D�g�TbO�T����D�uj1�����~n���������7v�l�WDR��m%M��
0i2�O@�p�vmz*M�?�_���Ġ��#�CX][�	���|?c}'�uE�ې>I�`r��gI���3{S���ʒ�yd�y�>�=Ȭ�|��q���K��D��������8 V J�LW�枵g�vD���q��hjtHѸEJ���V�[�Pz��8=��ǧZ�1%�����(4�����s���v����'�ҮAa_������qW��隤.2Z���i<�C��B � �c�pC��@�#�����'z��� ����ٝR"��'pt�Rj3l���
��
b����Do_g!�B�7�IW��#9'&/������[ؚ�ﴠK��>��w|jKsN(_�9\�[H+���V��4؀-����h�tRb��lU���P$j���h���c0�!k��{Sq�%��J��䟶_(�͆8(�奁���R��߀��p�A#H<'n;��*���ᖂZ����Uu(-;�'5��u�No���;��cG���U��V7��5J�fm��)P�Q������#(��*�;�D$8n����u�W�,w6�����>j����G(����ê����D&g��c?e�����u	�K�-�c�Н$gš�"���R7������gM��5��t&�X�z(H�=Y��^z���5�����|�P���_a�