XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+W�ߪ	�5:����W���B�Ta��s,�����Z4>�<8T'��@{[O����5�ks�ڋ�D>��x+],�ɡ,�&Y�#���ȿ8���`qw������'���+E��5#}V��{�����	c��˞��g�G.1�V&8@]�+�2�
|��	��v��Q�<�����e�jX%6p�̀T��2%
e���h�{�B(��/����gY6O7���%*���D�	��O�������wG�$���
�-��áB�Х���6��;��	��Ŵ����-�-̠i�Y�: �{�5wq�>�.�o����-cM@��Bht]�d#�ŉf�c~C:ݲ�	n���Q���x�2h/�V�#�zR�,b�O�2�¸;�{����M{U�yjz�p����0������ol3�YL#PXV��g,y�"��x����:��i�&<�8�g���T��|5�Ϝ�[�T��?���!�JZ���?YF�uo���a�tƤ��e��`�2ٲj{۪s:1l����1���PO@U8���tf��k bn���2���� T�m�⩨��b�@-mܧ|X�(���3$���\���a�K��'�@���p��ֽ* �$v�	Ro��W�������_�����=��������<�y$<T����Ũ�џ�q���$O�X�{d�MQ�x�_b������-M�O�4�wL��WJ%���R�%��b@���֠��k�Q�MXlxVHYEB    fa00    2030�
_�ƱDJ�g�xl3�q,�`���*W9j-n�J����A��� ����u�7#?����0�%[�ż\2N�q�ǡ��Ɲ��e0�ĩ�\��;>3,��r��e�b�@���dQؓ��P�]ac�zp�ZIߙEE�IҊ�v�$4�����@�tp���2�d
t��đd�g���ļ��ca�~ӥ�[���}G�O&��o1������'�Ej���ĉw�]ҥ�����@�K���d��[�ض� ����2S��Sw��Z��wj������)ä����q߆v� �F�; 5?*�Qz�/��]�	�Բ�i���s�k�$#03��L���l��E���C���~��TҶaE��,����-��9!B[K}xm�	h�\"�"c��.�-������
xL����s�k1b�f[��<sWK��24� ���&2�OY��ǿ���	H��YШ��<��8��X��5U��o҈W��Q���8�K����o �@e(g�_�,�_6O�%U���_�Ke��j�Qw;��.>��o8�^s�pGћ�2�k������u)�ݭ�]+^h��u
0fa'f7�!p~��/�-[��k�u����Zx�&9����@�X@��cy�a}�䂆b����0�~�sF^���<,��pn�p���%S����[����)}�)�?� �^{����;TS���/�Ȋ��*!)ǔ˛*�&{y��D�Z�z/ᢸҫ�l���3���h��/*��W������t�
��:Ժf�u�+7Bh�+-|�&uǩ?�|�L�5���6sz#F����,��Cc\7�>��hH�F@��1����}a��%k�C��o:7�_�ܦ��Wh�	���3x�bv/��*��a���ZN���OaYQ�R�'+K���ΐǩuH���pR'L��^�ǨO�="BL�-��FէZ��#��u�R<�~�k��>� ���`�+�~�kf�>�L�Ν[.�n���c���3˅a?z'���U�ü{|(ʣ���J3\c���+��0I)k��Xq"�����J�͂�p��:���Fj��D�&�LBx��i"���� ����S��x<3�4�I�´�ĆS�����n)s�G����d�X��H��"�@��������FA魭d�,,P�h02�%��H�/�<�� k�- �<貐�lC�|ɓ��V��'�%�||<r+P3���~u� ����&Z�3�y�햹0ź��8a�ۂ��b��,�J�Z��JQϩN�w��r}��,N�/�U<�g�,��	OJ��c�����3"O*�&��}i}�B�A�˱x��<�|�&L�q�-���ǩ^+Y����W[ �����J��'D븯۸���`��}`���I�X�(�zį���sO��0:�j)T��f���i�G�ȷ�i$���y���05ޞ����bCE��K�RpY�<@̨A�"�R4>�ԏ�o�W��zćo���.�Y�����5P��`~ �&����Ɋ(��r2��f�?�s�^y���l`��u�NW{G�}I�=�W���_�O�^>�2���B��Dd�1�����������\����m���߭9���E��	�N���ee0�.�L�\�7���xe����^�Ȋ?3�ہs�2�������|��g�tl@��B�L�";�i^+�_�}�UA��Ҁe3�T_�C�X���ii�d�ah ���F�\0�y�Z�d��ǉ��Q�(����K'����u;#{|c��$�-��3Na�u��$�����D�a�<6����(�������ȹs1����p��V��EJ��9�:�mo$H���!&tvN�u}��m�}��J��,g��s\��ҝ��+o�(Y� *}��m1��i���e5�Q��ĺ�[��$�"$�� &ە�F�n�E;�D�R�\H`e��E�����k�H��s6����W�xW�	M �!ư��=s��-8-B�]8��G-&ى���/F��p�e�
�ԇ�^ls8���1 ����:|�	��r��:� 1��i�+�9���%DH���5Rʲ�7�%$�"���XG�)�	V+����zm*H��@=�C�I1YGR�[�0
��m��b���ȍ�.-Ǿcv�R&���4ݿ��=%l�G���!_�K΁_`��=�7�r��4�*��Z�sB����Fꀵ~P]�����6\���=��h��Eގ���"7L�	���*e��2t����M�g����v��V{�:����8g��S�X�]sF����A�����;�!����Bo����R��\��;��&�V�����PR�_|���
��*>Q�V�IZb3�VP���L,��9��R��`�_D[��\݂�l ]������x;��������?۪�<Dn�nߗ0krN#�
G���g����ʐ2�;	�p��s�y�do����vPƾ[�>���0/uŰtƔ�|�rg�y�o�f�j*��0; ��ԪErDiEp�qv��]��9*��$�03���?{#9`�m ���|�Y�(s�����V�� d���ad*����^�G��,�g�h$��*���뚺=]�ӂ���R\��O�_�
�zт[�w9�W3��C�G{��� �Rlǿi��`?^OT��L�GfQ2��<�+�ư0ȶG�;^[>P;��\��u�KY�v΀����,r���G�Г>?NY�Wp�Z*u�����.̤����R�����7�p�Lu�룿��į���p|PT�R��}&V�z9���2S�4�JN���M�p����P�kXwk��i>�&�c�q��
�Z�FT��l��1��ìQ@u.W�E^��$6J�֦�lk�A��Lf��bO��&��/�6�D��x�˚f�KK@��Z����6E�Ԍ��[��d	��|��= �z����B�9�o�4�_������B㶌���)���LG�z���a ��0���r��1�^��X���&�ET��בZN>��F�.�'�|��\��y��b��p'@�jM
x��~P���fK�.��ڂ�YL�9{�]28���UH��nNV0��^��aZ��̟�|P�">��Y�r.ͧ7C��R֧��8V�V�����bo�T������:>����Oj	!�iS⦎	EML��	J�n<֒�~u}�M�V`���Ҳ���S�. �̣s(U��jU{�M�Z5�8=��LRm�
[��OlhG��[ �?̚B��	=��P##:��@�(쑵(���&����0C��o�р��Y�ղ?V�����Ǘ����U'>�l{��5��V��D
��D��3���|Hb<	;��n,D��6�>��e�!�6''��#���Z%��;�z��7����jѵ�2�9zhS�oҠߣ�W��88%K�i�B�ᾂ�Ks;�B���k��1/F����騆��i=��X�Ǧ�>�[2��d��c��F�~mED:�i*Hb�A��.5S_�� w��vG4k�B��dQQ&�SKؙ�G�C6S�2�|Cb!��T���Cڧ:�?|�CN�_A�rs��<�8PG%L��#ɪ��y��.u�h�p��*+� ��/'aO�I{�r^������¼�;�x3�́�wr��4��\�?-�Q�I�z�R�����������ҟB�l��e
���n��e"�@SL��~~f�3qf5�����'ۇr�IVW���\����܊�Q��x_��{ӳ�|�p�L\����L��(=���t��^^��F�j�g���G ��sX����=8Q�y;?><��W��)����������=��r��y
��ގ2�n ^����up�۹��y_$���1��;�R�߅E[q���_t�02Pv��0@�Fz�xj�qr�0��	���e��D��ؕ-UqK3��W��j�۱�_�,2M��,U��E3Ղ�.���?��u&�R��7�c���T&�N#Cn.��FH2}T\u\q/I�a޴:���O�(]�{t�,8��Ҩ���*�$,��8�����7%����FP��4�ŭ����#��-�R��WCSGʋWɽS ���Tb���8�)�E����Ö�'\�"��Z��/|@�"��H����(�"�B�OAw"7���,1.��\��I��1@-�,�@r��t��@Y���M���K�f���K/"����I'�~*�a��5"�o$�E�+�_I[��n�nU��jZmsW�>�9�k��5���wMs���9��D6t���{\��+���,����d���g�Ik,\����Gʸ.>s�+L5	��E�:�p'a��WP���D�������fj����.�!w� &�Ջ�j����Y�#��	�چWd3]I�3�F�:�������&�	c��0� w��P[4\�:�C)�|��g,w��izs�����eq�����b�hae{"�t'��?f�X��lW˔t>E����Z�kKK2�; eS�.����O�6��b7T�>���t�3)��!7�dm��������*l_�cm-I�[t;п��듺�Zˈ�1s�ǆ��:�siJ�p�E�u)�+=�|{\ǟI�W4[�f��ڐw����'4j^��޷��N#��ėD>�qēۀ^{tˉ ˘�O���5�=1=���p������[�I���E]�C���򌆹�N������]��K��8$n2�����\S����?Pˣ`<���(�KsB��k}@&ҽl��}+Ķ�x0�!��R3��-�v�=ۤ�%�Bc ϽI���׋Ļ^wФ�Qx>�]��w��~c�h���K�A�-���^����X��������x�!YEjA�q�j��B�f���u��i�'&�Pxړ-Z�9T3�I�OZ�rWf��G�)���W�����x��\Ҋ�"�����P�3��O��W���-��Um�ֆ��GS�
ݞ9�;���Y$3�eE#��ɜk�{x��\���,�*MX�֨[7<R:�!U,k�.+ ��4)���J�1}��x�J/�TnD@�U�����I�����$�p��(Sx5�z9W'��%�Qx��[W;��|}W2JE��z�a��Q+ŗmEQ�-��y�)Tkr4%r���	/7\5C֤a�q��2t�.�8��u�V�!�q�K�n�hLN��A���*��"RY�B�x���X��48:)ƱXX��Ɗ!,r��=�`Y�w	��lf�W�L�x���)t��kM���q�����q�d�Ҟq�Z����ܟ��)zvXM
����	�1�H`��3����#z�t������Dm�3�5����Һ����:_ݕ�4�D
��liX!>�
��Q����Iۊ{v(��pM�>r!,>��6�_�cKL����N���b'*]�x���C2[����؆!�0���Q���/�����k�B,��Z�
H��q+�BxzR��/Р)�Ĩ'���t����pk���s���(�z�נ�Ȱo ��W��������T/�R�_����h���q��Pd�ɍB���������DU�Ru��x�#b�S�Q`�|�v�e3W�]n2�F���hP�3���HD)f7�;��`
�mćJN¾��3i"z���2
�-q�U��v+ �Ubه�o���P�O�In�X�V�����	�������c�SvS�`���c}��{(O�X�kb#�( �!��
���5�C��K�b9n���^���3m�^R��R��B�`؀��v_�1��,dG�)|T�M�Y���S�e	w�^�<��sB�&о���ҫ���O�ځo(G;�j /CZ`+^7���%BNT�G�z��X� ����z="�G�WU����Ȋ���ǓQ�Љ��8��E���mjE8�Ýh���Xq@�*���er�˄u�ڱp`���
6��X��Kѽ����T=I ����1`>~��+�XҎS�
��N"F��S����(�u��~�-	.�Pmcv����L+N�������*Sd2�q����.��1����F� �/q�̟�Mf/�af3���@�M7�a-xj��O�a�����S+�Y�ȍ�E�������sͽ:H2��o��Y�^�_<�i�H�v���×f�|P'k��p�voTR��=U��� u�X�g�M2�w ����Y�X����l�����}~ӯ����������
����v����HA���-��2��䤋�q�z�(K������' �jxb��F�sU�^�q�!ӟ~ё��P�D��Ws]Z�o�~�9%},E��a�xs��GS���1I�{g;~{�N��,�M�{��M�-��2���h�bS���n��<�L����H'��~�"zz+n���^8��T��/�`�e��Sj�{�����y��%Bڼ% ǿ�uA���(P�]�Q���o��f����I�~%rH�-����I�8g�AY1a�4W4� 8�h:������  H��Σ�ԃtN�-����O���n�E�|2 y��n����t�kv;,b�8�,�yƶ��>�%�.�x.����>#�?�����m����Ҳ��6���^����7�U�u	Р�BK���f�Z�aU����BY��;Ն��[]+}�%GgL�BG�q�^���R�y�V�W�.V|ta�p��0�E���R��6�"�i��o<��9��!��f&"�i���ݧ��ԅ��2��CtK3��i�̃����ף~��p��rY$��WU�yr9����r����r�%�w���2�,�55k����$ꨶi{��^��+�7Z �e�w@��
-K�i���,3�M�щ~O���]k�KcI!�����KSH��g��7uhg��j<�z��JzDAc*��<eI�X5<ҵc�q{y�{�曞��Ѿ%ڒʑ���n�ԉ�Ƨ�,v�L$m5mA�ŋ�p�_xV�4d��JԐ$�vw���c�ϓ��r8���׳�=q1���o=�6$�/�UwJ&a��Z
���T;�D�o~���:�nП�o�p�o"���<k���L��Ju�����X���~��8� 8B� ��������Ng�$jWNIZ��֤7��:�7�Uܶ��-����q@��m�ۛ���]`�G�=��y��ş�hU��kDO��W
T��s�X��CZ�}�;���O�<��@w�K,7;\4hG�x�.����v2m����M�f,��lCph��ي4�B�Zp�7��c	l�L��x��}g�-�;���;��qZ�4T�ALD6�,>\I��֔�j�I����k���**>�X͢��N6�*ؙ�Q7Tj����&��HV��<�p����K+:`'�7Z�G2�{��(e�ۡ�6���6u����#��qA��c��fTCʰ ��6x�NP�`�2��1S�	��P�6��^�X���{|�TA	����D(��
txE\z�H�YD��8����C��O��� ��Om�y��dm��V�]6�������1r�TZ�)�ΰ8[D�uE��Q�E�_q�j��_	f�Ј��1:�t4d�p-�P�qP4Z���y����!H��D�"�T�T�RŉT�`��Z(h, ��T��mh��lq݋�<���w�܆uG�p���2{�6Z�9���_���8"&[5R�7���6�#Ofu�<s��zS*8'S�.i�����!��ѓW&`x�/��
'2���){⢵7��e�$?^	`>�ǟ;���T�-wk���"�������Ш��Ѐ�I����˯���������1kwSt&ޅˑ��Y�J1�����a(>e��Aa�q���%��EV{�����A!��)8Z��?*'��00�L�xR�gl��=%�YF,�Xˮ�۹��N ��q㢒��w"��Q?״�œ�qe"��2r�*R�Nʖ=��]A+!d�d��-��ڐ-0�U��?�i��ф$K>�d��sB���O%��m�5�����/�H�������6��ܑ@�	�<���������z���I�d�?�r����5'�� ?p�����v`�\y�t_LM�'�������Y�+�x-L�K�y=� ��4��s��u������*�]�XlxVHYEB    9620     d701��������׉��]/)�k��Ʃ���r�x��k�u��0�ȕ�b�Eɲzr�ʵ_��1�ۢ��g���������*�8ø~I��Sm
����}�0Y�TM�q�5�,Ǡ8�蝧�N8�ݤ�kO�.�睻�o	a��j�8�,`���ŕ`�x����u�,����D����F�]���5�������R"�l
F�
FO_�8�ݯ����6)���#)Ժ*װ�:9<Y�)��#]f��!:��A��	H��y��wOr�IQ[_��T���a����0	8�5�x����-F�K�Z��6Q`���]�x�#�^v\�;��m�Rih$Ц�j$�G�֕3Z�ER[�^�	�7H�4-�&��b�x4U�;6@�Xt��LKTʟՠu�D�ǣX/�M
�E0�&�nV���S%y{y�%$/�跒wμ󭎧�+����.ip�F���Ԟ��
�Vᚚ�b@z�+�C0�MR��x�Í�$�`)ڬ�'`]�N_�X�c�$���D�л--�@o(�V� 9�#?��nՊ$_�N~~'��hñ6��YΌB�۝�ip�~O�.�������0��3�x����H�W�fw��m���y��w~Bfk�<�����m���u�ǅ���A:O�G�=`:��5�����9�z6+��<�V�2��و�t�&�+G5Ŭm�$LK�g"ņ{��ꩈ��h�y����X���I6g�Kӟ�P����gߡ@�K���z7�V�4ȁj�1K�P4;�6���h�"�0C��RD�g�A	��y/>	��"ٜs�2���I��]����	������zA"�����Q��9yć�;��Y�MIw~�u�r��B��I}�d�Gc:�&�&1ݓ���B�9����L�l�5���֮%Z!����ډ�Wˈ%M�T�q����>��a��u���,��q1 ��]�a��Ӥ�o@�(�G�D	���(��.���f5FK8�0��մA�[i����OR����ceZfR�ص~h��L�X��Y֌���a�ಽ�"S?mkn�E��[ʁӦ��N�?ޕ9���+�
�v@��s�"d����o�G�FC���ZYcʚ�6�U�j�$&ζ�p�Ѹu2�G(`�*E'E bn�}�D,�ן`�筦$'&�yRY`��ix���V�;)�qG�?F�Hl1����ﮦ�P������I�ic'�t��,>∄�"V���&	�-fn�2 ���R�u��"0��@K�p�6t��b8�J7���
�cd}����_�b���T�0����m/���1�xA֑X3�+v촦���e��\�Hhw��QxyB�G�"�߱�� g�8���_Cňg�57BU�g���uay 2�5{'E;�+u�&�p\�r� ��������wB|w�Zս�@�(�~B=�#a.{W��q�;�c���[-Q�8�? �h����� �Z�d^ˍ��鍚�ҍ��n"�{�)�o���9nOhĜDD�k��~�ҧϫE��,Qo����ZEYN�cM?#�yP�?���,��[�	�g9�טo��ϭ?r���$!Ct�:��On`;����AN�bK{ٸL��ƔT�v�@��
��GZ�ς�Y��Eco��y�)�}Ѱ�^R	UU2+G6%�V�L�9%�v=xᘞ�'�F̽�k`��Y�Ck����H:t����B�T_i[��D�D�_ ��,3dҢ����7�-i�Ҽa�Մq��Cz.�a���u�&�"�X�?��|�0?|G�'�ep2��[�$�v��i�.�wl�B��S~���3pֈ�|��Ak���-�c�W�s�����;Pwq�\oS��}6I�<M�z�m���|���S�S�6,������#Aa����ZF9wvy����H0&r
��7Wmx���#nOi垴�ރ�����k����lrG��R�����\��5���鮱�[���ѿ~��<�
��k �s�X��i�4�4:h���I���<�Nݴ����v�Xq�,�ʪDӖE.��?�}%�}��ɃI|x��S��`�k7��Z�@�9q8$��et����W�pA	/h[o�~�@X���A���r��{��)�a��L��:lg�?�����G*lw���Y��mD�4T�]Jg~�]ߝ�5�TS㾝���oa{SݑV[�U�YN�t��h����>ʎ�n�@A����!/2��[Ä���R�AB�A>�p},;f8G��7�ׇa���󸺢o���W�d��8`�����O�9�g
���ԴĞ˼�y����G=��R`�1�R���Ce*Q�x�x�c���3���:Y������C
�i�<	=2�8H�h�h	�I��mc�1:�G�dW��J��-!Tr�
��CO�hg�?�~�Q�7̇��P�넗�>L��+4a��UT�}䶑!\Rv�<b=^�Z��nDќ)����o�M��̲�j��-��_?ckJB��� �Pj�b��b�r��'߹���W�"���B��q���k�͉��R�(lS��i/[\X�8��X�w����o7���9k�;lm�bY��v/�v��[��Q0�w�)&����^C��d��05�D�ʇ�� ����oa�y �����y��c��h¸�봽�Yc�����4/6[��?�W���q1^���A�1'2ˡ��^ d\aDSU���>��zjRD�\o2k��f�sK���F���E�)_�?�����LC��?�|"��Y8��|D����/״��Ǣiɷ� �2�N"Q�!��Пk?D�����@�*���j-�y_�`F|�����[��.}�u'\����,'����i׼H�ګ4y�+��	IT�Os�c���{�|��Zuߵ����4�����|N5f�"='�N���K���]&-�KZ�cc�:{U�򛰃5z� �D�Ҽ��x��T�bK�OX>�f����!2������\�
�lTX����R���s<.��4YP@W��;T��u����s�*p��=\������@(EB����T*�h7#a
��e(��趇��Ѣ:�e�W@}KP���R��ٲz�dD�Zw ��-��&;|s���L�T��.��_0���l3���,$	��O�W�̉���<��4 �C�����Z�L�+/c��>7�D�����d�X<���6�1��1��xĀ�}Ƚ���G�L�(�܀�q�&�=T���> st�px��P�p6������&J��s5(�XCdc���8����(�*%=L�'�7b��? wB\������l�ڭur\�.�02��v~�EW'�yQ��@�
y�Ƅ�����Խb��Ip��N2i�Ց�@�zXi��(��!\��y!'�����e@iOP����e�"�{�6X�Ei;%.0wQ��=�Ȱ���Q��