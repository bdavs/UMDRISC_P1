XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���|�Ib9��T s�0�ߑ+>z�k��y����moY2`�;�/ڿS8U��%�bU��(�G��q1(�2��@Q����!�f�	�:�U�[� �SG�*�4-�qgvW��i(;���UUvm�,��.g�cWu��b���=�0�~�����!Q���c�ËD���=��(q��q��e��	��]���0D8�y!��d�eu��Q�瀟o������R�|˲�DU�YX�ܸ�	)_�e��.7J/!�E��������,:���_j>�}���l f��l�Dd�����[������pw$D��jZ�<�t���<z?Yئ|�� ���P�ax:�F<	0���H1E ����y�p��)l�W��-�KF�>�ve� Iss���ɀ�3*��FY�ބ�&��]�-�ڙ�&�h����" ����3-�F��M�9�����S`��)�0 2��w�qXɝNÒ�3�I�����(/�O#� u��������HA>�&���(����Cr�/�&T��1��s�g��#Q�o�L�az��(yK;4x�S�2
QȊaI"���u�,�
���BX�
/{����b�l"2��1�i�E ��.����?Q�"�@�yeYK��^6{=���rmS`������o���a�R�����<k��^��b�p\v��9o�=��N��w�q�rk��F�hۏ�4���]�f�`����z���X.'������/���Me������t�]�앺!\n롕g��q/-|9�0 ���sXlxVHYEB    fa00    1ca0.:Û��lB��z=����1��=���fO�֔�I�HOU��ۦr��!Bss1W1Q��Aq|Ap`�3�����^�0��
4�b�e�F�-�Z��ɝ2�����`��+]ıH��Ǟ�Ǽ 
5v����x4�I�r�ef!��S ��s!m�u�R	;���v�.�k�j�v�/p��ȣQ�%E�������'�g,�C��,Xxˢ�+���Tœ\8���ϟ��Bgc\���A��t:�x��X����]{J���p���xD��Z"٪��fg�D������(zE`�L�0�k�����?��~)�ϖ�a!;<�:D���U�(��S+X�f��u��X&��A(e��c�=.�0�je�g�����Nu�ر�)��%J�S#��5���ً��XY:�	��9_V�����O�T�TTkӼpk�l���=! ����%K���F������a�AM�� ��d��T�����-il
�Z����F��I���T�imI[#�uskO��в.�5�� ٘Ǔg`ITM�u�T��V���)��i��tQ�JHj�����{W>BoY���QaԹ��I����_�;��mE5�Ԕ��N*$�'����g���=�Y�z�k"ʳEVL�(���UO!��5b��ذsr8�x���a
nB�ޛ@�! v��]��A�/���ዚ&�'_�:3Є|��=��dzBx�R���EN_�}h�
/���}�^ �[g��e(�%V��]i���JbX;=@L ��U����xk�@�u�e�\&
�8�*��2������B��V�[<���̈́�!'P���ei��@
󣤤�m�.9=���Զ�i�E��ʏs�� ��$��Xɻ� !�j��.�T!H��L�&k�^Q�!v,p.���2#ĭQ��8���f��(��g(Mr�w>�)kdl>[9�kD��;s��^��$9�W�6��$<lHڅ�JM���L�&�܉���"�g�w�b�I��CsIf�{�I)(�o�Zj'R5	#�������C��� ��G�<��9^���o?WF��~3�m���E�vTO�+9t߇y�oZ���ǧ�.1Sń�l ��#�p��S�wC(���hX�P��.kqb��D�����?OQ4�.�Z���5��jJ���Zۗt�1e�����Ʋ��D	�PE�+=�[�� ����7�9_Jֱ�[%!�Ѓɫ�;e���ph^��>|_�4B��H
��&�HV��}�Ε���%��vR܅֑=��GM��.f��a?%=�Fs�]Q�����v��/��cUL����BGv�c�ǽ����ڽ<6xF�}�<q���3?�ǢNk��ʟ���d����+����X��o����U6+�T���=���I��m�]
ӋB��.�rV��񬼖_e1�qF�2�B�Ԓ7h:�@��3�k�8�n}�;F���K8�:$5M�d�J��A�z������������M/?Hvz�i�IF����$�����B0��B����zqRG�M5��A�)�\jO�V�G�6B�����n�4¤zJ{����Xz�i�k��<���w�/���Z�V�ҸwhZ�+#�����Y�K���iA��7�3b<goY�|ʮ���h�yBO�?&ؤm���m��e! jp��`�g����MX+	r�wBوl�Zݑ�<�l
m�&����4QCd�Ҕo���5HV뱵����]�@�GHy�a�@�'tGd���<!G�d^���ǋ�#�{�(�I��+L�*3�,����6iֿ�	¤������m�����9V��H�,�>�5�,��gC����At��V�S{3�K������S�{��\�ߊ��C���l�W��`�"3�7h,�.�J�l��9F!@�Dl�W�H���^�M�b!Fo�W��T%n���w!�&/����| ����5�����l����i����N� �x�5SL���wq>�p}-;ے���eG�;_j�� u'�w��(a�"4�͚�T�f8F������=�Hhlx��k��f6'�E�.���&��fi�����(��5t��n��~G2K8_@�fk�5���*N�9��ޖ�ёMP]�*=�-���� |�]ͥ�+l�&��`��$����i�Ȭ����Q�~ס����n���k�L�O/7/@���i�]\/:8��NۋDc��e�;4فcA�-*S�ㄜ������I�.T����܌�Tq�V���4�R��$�Nv=4�BS��D�wD
݆E�@Iɝ��Ug��M�g ��Jc��<�Uw������3�p�e�ƙ�fq���@�#����R�h{h%�_��?!�?z�M�����DJ���.�M�B��`���jj"����@�r@�s���.:�W�r'`du��o~���6l�1V~B � ��A?V�)�3/�-��CU,��Q�(E+����o`E��(w���_��ZL�u�s�ty-B==n�� �}��|'�.^[x � d#nej��&�FGT퉬���{��[�)�������<~�g���2�Únwg�7s�)����D�
~=/���)�������=a��[׮�]���^2�� ��<Me�{�[Ȕs�d!|�MtH�? Y��dG��}['vfg��B�݁[vm�Ό ��b��BF���s��.zݬ�Ox���uf<�7hJ{�n�{-%a��q��,�2w�@*�AV뒻�&1!{/��i�g/�Dg8�"oHdY��D��\���@��qۘ��(9f`��~����C7�.*f�P�eQ���찒~�q� �G)pT�y��wO�śI��#���[[�P�A�7C]����ʟ�L���(�����v�����1�F��q��}�7!;x�D3��i��y�5�g=��ۯ�#U擶�}ΰ�p.��Iq[Z��;�;I�pYd
z-hK&�1�M��Ռ� T�5O�Ԥ#v!�����v�_; ��%7"�<p�h�0��}���>��ޅ�&�G~����Ԁ���"�Q,�Jsȱe�h�L+cj"q��cd� �e>79K�Wv`���1�y]�i�\�_u�;�P���x�ϳ��Z��vS��v}K�'���/L�j�͢���n��\!���f�� �\�Tjd��se	ֺ��C;l|�hf�Q�<Kㄏ!	�"��|С���XcW�&uO����p��ؠ��P�Z�( ԋ�G���6a߄�KA"����מd��UȬ�(Bs�D{�T���M�;Ca�P��LiH.�<�������V�O��B���K�@���d��o ��TL]�4��8p���Wh.l����6�!�'�z��V�i�rT��O�i�E���^~�-�/>Kyy�p>��*�re�����3Yy����~�ٙ���
��>4rh�x�����qG����F�JW������1�ţ-G��<�H�#:��g�ai�}�g�R~x��#�[9�LK�{��Ta��.�B�7�R��罙�&�qT��s �1��$�g@�j`?�*V�,Ar�e��#��^겵&���5�B�.l3S��(ůKuD̶?\{D����8�ZϘ�mM;,Ϛ�ن��eZv@ݫ�۲$YoA�Pcmf�T��mQ�n���d��^�.)�ey��˂,���=IY����x��Fx�S���a��Ww�Υ�b�M ٬���{�	�Q}v[AǑX��R�h�,�v"A�d�	݉���2X��� "U�.�3�g�[�^2A<$�7s��ئ����~]�T5	=�x�G����XwR1'��UMRJ��;"�dنxc@�:�6�`�*�����K��^�{�NY ʶ�LY�A���<-�iGOm*Dđ�MU8W�	�ha�ߥy�q*�q�3QD�	,{\��� 쫢S�?d�Y~ȗ��o�I*`��#WGЩ�d���)��N��[�8i����m��+3v8�ĳd 5��1Ӓ�O��PqD�\��sg��*��n��p�r����P��)b��dS������چt:�֚��dȅ�g�S)��!�+�=A�N�R�jUCT��T��d�x73�B>ֺsuz6}#�S�-"u_�$Q���]�w�l�c*x�� =���Y�A0X��Z���{���˄�QK�N�3ZW����G������,<]���D��b�v1
�.���6 Ď8�ɢ2�2I��
8;̇��Z:���>6*�X,�>��'�l��F�嵻��-	��by޼|Q�ƍ�U�^9'�P����0�ӈ43#N����6�����B&
-���y���W�,烳̌R�{8�SO���	OT�r
���*s����w����=�J:��U17�{���Vj�k�Xʮ�D��/���?�h�,\�&�w�P�Y���)c:q?U9r�2Q����VF���s����k4�G9pіɕ������r�XL�����˒"�f��3OxWV��5�tǓ�%�5FL׎�l8゛���n�a�:ନ�j
���ԡ]���a��8�u]��?_�OH���ƈ����ݠ� ��{�7�_�AR����e�:���f':h@��h���Q������-�=׀}iY�5�����������,�V�]n��=Pp*�G���l���0�9'�a�[�t�yTWI'(I�BI��3�1��pj"�V����%Vi�#��P�tp8����n���&FMn��4���8lG�+�v����^��_��[޼cɍ:��)��S+�f-�eݣ����>��À?�g���8ꔷH9�I�>+-��'0���ĝrƽF���8%��B����!
B�P����#'tG�TR��	oܪC�"T\���|�׻9��O�G�
��9t��Ƞ2����˘��.n�LhE���*����Z  X�Qo/�fJ��д CdO����'I`A��I�?�(L�K��Fw��e��l
'¼.��b��T��tӔdg:5m���2=@
c[|�A9ǖ��3�`���&�:U�0po4��
�H1�ָ�Jbe�ݦ���v��RKi�ٌ��,�'}�fVgP���tC�MB��j������A2�&�/Ka9�M��!�=*z-����^��L/`��T�MV�[��&��ľ��|�5�tk���k�C&t�<`�B���yy��L���I��P��쳂�g �K��({s3�C�;�S�hX����#o��Y���Zhޚ��L1)��m���C冭�s~hęҶ)�%�%b_	ԡ�)u���>���>X��h�d�ӱ;��J�U�)ީ���	��=8�ɪ�ю3��}��"�9:��3�_SC��z��#���$jG5�[C��ڥ�8�={,ܒ ��D�{�b"6�J`Z��b��
�>_��ղ័Z�KXu��ޠt���!�@Gf�n��o@$+�*��G0�x.o�U���P��1�����P?�U�R�B1+D0x�(D:P�h�����GF#�ǲ�`��Y��ֽ�Nƶ�5}.�m��$۠�d�[
p����7�*0�c���U�x;i ~�
Z(zwKGoi/�F-*{�Y�Rm�.11�XN2 ����I 'ц�ea�lx-��G����$��|�M�M<~�L�����]
��s�s�@K]���S���F{O{j�SJ��4��v_a��ۼ@I	+��[{2������������/y���c�x�['c]>wmو)%�\<�/�ϒq�a ZYC������:�խ��l�V�]X��sd9�L�h0D�9�]������zo�y1�P,8tH��~L����	
7y P�jAb�B4b8�'av�hW���$u���������� &ܞ�ٹ�O�5�<���)�v'�Ϭ��� ɏJ�o�;�͖�(�1�����t��N*%Cd���S��x7��}�8x�[�:�&�/��2���S���|%f����ş�Ydc�JC�2?OF}�5e!WF:�pUi`��K�Z��ޫ��i��O�.R��n�x��.-Vxس�tڵ97��:*�B7�E��Й��y�x���O���7��*Z�x�����i}7�7��{�\�_[�[5d\\n(�P,ࢊp�P��Gޕ��y/�׀���P�C�X��#W/�c���~����_��:w����/s,���?)2C��e�XK�_P�W�u����9�N��붵�}�]D]�F[�mN�G�}j�_>�s'��S���
ƽ�/�?� Ua�ٗPj�M��k5�!��y�ט±���,A�<��Ф��W��ï������=FZ#M��8{NJy����9��<���z���>Nf�	�XpY�B42��_#CP�?"E+�Ȃ��J ��o}A̓�36�}�c�P#NTܾ�[�稂�_1��H?�m
`oi�]ik_^�f�2���?��;������W��JН��g�Iި��*@��o?��3L�H���,�^�x(�HY�C�Sp����S���n��a0��Wz���
6bרчa�~f�m�%�l�]�<3h��������#
@g��%��d����5!�7���ÜW6m��|�&'�k��ts��!^O�X	�{��(��d�uh�C��M��5��[`�<�Ҕ��*K��*hG}F��������|�������p�+ȚJL���Ny�L�Q�w�Z�S��ᵺ"�F~/Ýl�7�X �㙮�%��y��5�Ф�/�G���cݏ��I��Bky�㶅�Gw7K)$�]s�_�*�$�ơ�����6�q�� !�dI��G���A����/��}�P})Y] �L|�D;��,��l"���!��w���tP���˧j�r�gF�b��U��-��l�p����{,���{r���zkEj2|��������r8��ƈlW���-	���j=[����3� ��t�)zG+���P����%�_E��t�,�fvB;I���ܢ��&�)<==M�t�z�)�#lƊ�=�5koU�@�v��k���wX���=n4����1I���a|ݛ��lyҴ��ÚO@M	�~?7�������(�˻6_ �#�a����t�����N��r���<�#�kt�{��k�B6�4k�]�˰�\e���3^!����WJ;�=sTOz�K�:B/W�\��,w�EJ) ��%㐹�
;3�'�fW\�-)%�oy:n~A<��DG�P�d��c{��XlxVHYEB    fa00     cf0�e��E�_��H�0��h;��[�����Aɏ�˻iZ'���6i����۵�k�A���`�
\���M{_�2�� !_�:|q���^�;��J{oq�vu�D�UH7"�i���b��E�;�@�PZ��$�kWIڏ4�9��lI�s���դ�:}��*ǟ��h��f�=��9������FK��,�-�
$a �npt0S �h\Nl9�Ca�>J���>e�%�>�wZ����N:Τ�	䱋��p,�09E׻���t�6��Lߨ�ݑJJv��90oW-y^/T�v=�flH�wl	Oŝ�E	�1C�WQ�v@���7��X@p��NJΜ�ݛ��'�SJg�|�#=�p��ʸ����X���ǶxN�� �����axp�*~��Ƕ$���ŎH�2��͇�"x�!��C��K��f68�e?��dPfd�=��[&�π�~s��yv�u�����͝���)�FnH�}�	����Y��E��ь^�ڐh��XC��
���;��`V�j�~�_P��@|�k��Yv�F0��H!�<Q��p���8z͑�~��)�M�����5����q��ʁ�k#�"�m@���.�Ʈ��W~�:����qm+R9��Ҭ)�ςX_����!����4ȓ�6v��B������Ghl�;5h�1��PW���ktQ��NuWQ�A�_���q�d7`�� �WK���{gAȃ��8~Qּo����%�"��鉶 ��4�֒��Y4�DeO%�&Z����m���@�Ű0D-ލ��2��i,:���6�H���35i�z$�zR���u��LuRN=��+sI�,�_!��C�3|3�B��������W��������1-�/�C|�"����=ک�w����S5C�4- ����C�'!���	��P4C�`�C|B�F�n�����}�Y�#������3�v�f���s�y�pj ��|�G�8�(BÄ�܋&����qZ������M��u������(�	�hþ�z��k�?u�	��=i�+������{��	��o+� ��Ar���`�s�)�Р���(>앙s
��!{�1�"y�3^_�N�b�٩�;X/�y��n����k�a���k�kzwV�?9�,}��u�ap�W��y5������-�� l1k�]�K>��7�|�(��l��3�#�P�_����kz�q�^&)�����g|����
�zg�(�U- �@������N�6�5����5��ٞ@is����S�J�-w�h98j/��RP���:3�:B�# �/���t8�����h��AȀ��u�z�A�1ܴ(�5ׅ{��c�q�����Ů��C)tW��Łн!���S�H��}/;��f��m$�a 6Fs";3�o悻aqej�tH�$�3��-'��D6z�:HNBs��qh��#�dl�L��
���Jt���j�Ҳ��G����d��Hl�Q�c����R�5���C;W3�"�j�2�w\���Ƕ�7_>@o!�:�[����Hc�]ê��ı�DWE?)��	>~�Q�t]C�q<�����Y�
o	��[�f.ɠ�õ;�Ó�	N�ジ>�u�8F'B<ЪӫH�L��@O0�;Dj�wm�a	ʵ����BO>��)�4� � e��E���V�-+�a��t�x������|ס>k����,�
	Q�uW �����g�a�~�)���M|��A���Kt����d�two���e��QpP	#�ŗ��_�#V�=OBa����1q�_����[�����?r��4��v�B�U��Gy���0��`�E,=9���m�.2��A""��NFI+�4��vX��Y�����_�F���g`}�+Gf�[�a�`�Q˨=�*J'@�g�aJcQ�1W�b�����M��ٷRPe�D�#��3��P�	m�-�7������P�]����e�3P�C�����Ni�)];�h�����[v�������f�5�fַ9��e�ܰ��>��+�n�>3.3f+�J�:ݛ�����Ajb�	n�~�/�+?LέL�\}<런��	�O���w��Z���V�X��I+�K� ���(t��yN:�0Q����Lk��4�J�Y��Q!�I�;����(�L�n�}%�")`�+�	R�}�� ��V�i}yPmԆ��"��!M��e�}�ʐ�� ��!d�a	Uv�V�-l�L8����6P�8G�<�p��R��6�늛�0����^o"1z�����U��2�ݾf��;?[a�i܀��$�萐v�Q����R� �rz�%Ys�� �����_Y-=�%���o$�
�[K1�1�w�s۝� [0�uk<x�߻��'g��>X��e�[e5sn�_BQ�3M���q-7��f:�UͺD@4Zn��_��3�ގ$] y������<VQ�5����a`�!/nC��@Uw�KrQx�Έh>RHn�)q�I7e���­��Y�~�R� �%���d##�N��U�o�N�^�X�T�O'x����T��+j���x�fo��P`�T=!�F��V/�@�X����ۨ/���Ͷ�g<��$���f_?ʥ�¨i?��� �@Be�#}v/�Մ��0ܖ� �&�w�� �R�iC̣y����Z�����������D�ˬ�8"�3'�J�x���(k��p�hav���A�dӼ�E%LP
t�)�,�@/ѡt��vS ��������_��E3@�Vl(k��5m}94WZv�l~�[��*	�);�>������ Ԉ�8���]��y{��q-@3/����lp�l�t�_�'oCTo20OIod��/�>R�s�lC��������TXB]RL� ��G���Ӽ��(������ę~�!��R�1p%��"F����ط0|6���p������&���|qw�o��*4G�r:6"_�R���SF�n���������g�o%/B�o���WFԥW8��̲?%��S^��`�5|���P�k��8Ut�����;����_�X��[ ��.ba���5������3VPJ��="���H���hq���8��✨���P�5x���K�hdD.3�~McU�����V
\�� n���3��\s�(�z��;e�J��2�j�q��R�ѣ�WVl�;6����+M�(��𹿮�����'H��1ҧi�U�1$��ZO��q�Ȋ�m�x$�ʛ�y�8� �X���Z����T�3��f�12n>1B��%�H$XlxVHYEB    3981     4d0'�)�R�5����!A������Q2�P��{.���7 ����Ǔ�I�	S��1ጻg�os~z?����kIx�%CE=�\HםEbo��������G�w#��������<�CM�XP��J�ؗ)�G#�kͱ�/��(̷�,�SG�\��<V*��/��BpMTӑ`��ۄ�O= �v7�xn���<@S�J�F�~��R�3{R<v}��J�rJ��H�9YGx�0kRÚ��|�|���)��
N�qveMC`��`�����	c3Gbl��}鎳�H�f����ھb��o��o�Q"%���:a� d����3��1��v�^2�M���錒j���̢߯�2��~��'u��
�ƚs��9�Cq�
��2���F�0Q{J�&���q��$�m?����qQ�&�HYG�1�d-��� 2�&�sH�m���N�Ćғ�GMRFk`Ɣ�o��ViW��ۮ�Î�V�5�b'�-v�v���0�$ؓ�]��j����1�q��_��T� |v���>�Hw����ëe=�f���V<0b�p��Sa�������,P�Dki���T�j݉�`��^#;��'��\UH.�%�&�<�D1z�(��`h6��8��p�*5���u@�,�[֕�ձΆ͎�U7#�����n�ԍ�d��]���/�bpaE8�Z��}ܑ�F g��z��	˗݅U~���io�$d2P�5�@�+����S�{�w��X�SI���m����sh)���U�J�{U��m�����	�=�E���ĩ�������Iă_��7��t!�Ի�8NξU�O����Py�?�1�7�.��J�Y�s�7�ȴ�"R���M��j�%%�����,&"	"ýd�bY��%.�R���=f����S6j͒�+�&�u҆�F��G��H�&�dGVǣ���n��;Nc�j�*��X�����X��~���)i?me�i�OL�ZϘ�ء򫴱�h4�䪑B	�5�! �����0]�.��t�����*�c��VKS+>���i�j6Ў}�qX�yOZ%*Ї�j���X����Hѣ��E����e���K�tf+n�ز�:%n�!+�XOqy�K��6Ҹ�ŶH��1ã��SlE�0�n��,6r����aV�C9s�3�p	|�q��s�z'�7"���J���:���Г��} $��J6T�8Yմ�$����O$>/�_���