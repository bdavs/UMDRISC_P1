XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o^<��VA���˅��o�p Z*��9|�^�a��!�@�5�Q����ZC�5�� ]�ګ�}�O&�^��X'��eݍ�@�Z:����֕H�<���C�6��<Uc&x��*-4��>��u�og͓<��~�V��|I�0��Ƀ'��l��u[K �]�+����s$�`��tLm�})`c��i��GH>�m��Q5"����ǀ3+ B՗�z�C�G���&I5��;��D�V뢀Ȼ#-�ÛV*�~��0�_F�
P�24[�Ʋ�ȧ�ulU��`��� �k���
�G�|�Zm\a�`�+Q�p<�8��sT%���3�!*YV�:�-��zlx�jM9���_o�q��������n�ҷ��],���_�������=g@J{MD�;�����DL�b�|�-��߁���M��Z�n?��|F�
���}�1Y6�i jM�p��D����J
~�)s��h<�D�����k�$�S����k_b>+���y#�wvۃ�A�aw���#����n��\�$��V�YM2LU�w:������g���;��`�ʭ�&ޅ��"���|��y�2����a9��h^����Gu5�{���l�^C�R>ThJ�Eߥ�X��s�3]=�& (N(�X����]�k�ف1_�q\�Y�~ax��o��8N��,8��WwH�����wM������%�&�t6s6�*�f������l�疚�Q�}47��.��9>�ٌ��6��g�(^��o,t�R҄��XlxVHYEB    fa00    2260����;5�i��M�@�$�Z# Y�b��*��hH6����F"(���/e� �'%�=��}��	j$��1Չd�#��`E��z߁���3�F�j� '�.[�Px�[ɤ౐A��f�[̇�Ԫ�9�"2]�V�ꁍ����y0H6ǁK���2�D��yМ]���p#����6�m��C���0L�s��yivԂX�"�5�EX�O�Lֱ���4�Ks��%c"��[`\��'�,����|�.�o(�x�6��*���<��;��[�8L�dȤ|��
1���Q�xh3e���Vy~��j��C��V��ʇ4-�==�@���	��?���]�����֥GN#b�Aj�b~�o���ey� ��|���:kE���R�������Rs&K�b/�ȡ%u��yO�u�,�"���Fp��QCr�.�{Q�MQ�'��8
���uJ�>��L z.�j�u[.��h���$�:��B���q�>��/AS������;_�.(Z5�3P�+1��y�tm�:�3��jƇ��(h"��Z\��.��s .c$͌P�=H�h���ȉ�_�\�'��{�_y|��~� ���ټLMg��d��6�ݎk6+| ��b�&4�4�]ORhV�!s�������je�+n���]B���dߔ[ �!�b��En��<�=5>Dk�|�݁�j_T����ϵ��pI8YD�#�j׫���w��E� �z�X�������6���-o�f}��KS"��H��>���k�[V	�w0 �XM}��1@�
�g`���n��%umИ�'�����P�|C��?���b�,��3^?��@`�J<W��gk%[� �FS=��/=�E��Ғ�r� �g����?l�T�Z���V܎9�F�-����'L�8�ԕ�^�4:�9Aܬ�Y�5�֖��ؒq8���1�D6x�I��� �26Š=���x[K�>���`�x�_�A���� �Ih�.;�P��]�&�0+�<��	�F�ڋt�E_�8f��Df&3�_�+��|-E�,žtn9n�+ ����lD4�N�~~����E .Id�`&c:c��{��c�������ᕖxm0YoS���Qg6,LU g]��KN�����|ƍ|ȣ��bi����z.�m��d�7�,Q�d=�].�l�|�! |��Bvt@#^��*��I�N&���Γ�xy�	��b��O����'�[u�v�ۆ���-�����T�G������A%͈��x?(�����3su8ieP�K�����8)�qr4F�#nU`������4*�A���9i���d�O�Ҡ�d�V���8�t�΄�����sy`LX��;���@�٫�b��a�����̽����kBؿ*\|ݘ�w��D��O㰽)���ɘ?�ͨ�b�4487EaB$9]�fIۯJ�T�\����F�� :�����'8�nuj��[|![��Ve��&�:�FzQ@I�٣��HaMY�����1w��u�;qq2��RЮ�߱N ���C�$#u�w�ZT��i|� ������E�� <C��*(7�Y `��ڗ,鐦�zs��M���@��4��`, ח��L���|�jF.kw�I�~��7��8a�J u��+��䱉*��l�\y��<܄���L��	<�04�BU����nq;�ؑ�x���dWs�%`x��~�>�uR���Z���Ю#�v7Bv��J�W�Y,0�~��Aޗ�z��8��So��=�{��
Y�OE�f8�}���A ���o��E,O�Id�`�7?vJ��8$�p�\#��O��:�K>|��d��Acڝ: �1]2��Ohf�~�̊����11��l�6��g���`�!�����@���(=�����𹦩�]�В
�\(>�ȿ�@�gZwݗ����v{���*ϰ@��;�\w�� _qnP1���c�^�7}�l��n�ol�l�ϊ����.{d����/���^$�[v��E��;�6��5��y�xD`�%�N����?FD8�no�E0uT���*hm�7܈��-��C�H�Q��:����j
�5!Me��=�d8A�ύ�4���8/v W���L��/�����'�S:|�`��cp��+����+��WZ�%��DϪ���w`®N �u�T�F��?EsP��X�]��/��Ȧ>�m���|�T��n��=�A4�2	�䋭b�Q� �0�|A3� ?��wT�s�@<����P#m��)��
l�KexH;���l��%�w����f��b������cP�-�<d�#�XmU��;�!򔡺��m��p��
p�qi�;�b�;��h��ρ>p$ȃ��/�)��7JG���LM�a~VZ����cwL��	���*>'�5�s�W�{'@��t��k�;��>��kcz|Je5�'����tk�x�L(ztk�>S�[D�Ќs��:�_�x�1[�����1G\�K�I�?�L�
Z�/���e��	�eSe����n�j��C�A5&�@�|�u�����C� Y;�P�Y�,��
xݸ�{IG�M�H����$}�������ᅵؗXsF'�ve\>�љXI��o� }����':��*���g�2�?JQS�
����/�l*FRwa �fJ�D��#{Ō�=g������J��rL������a�C{�n�#>@!����O�]���A�;���
�E��'��yM��5=��7��^"Ρ\Wλ9HјJe��Vʶ�.+f4񦌓��z�{�-�#�]B����m�mE��s�x���o�B5l�Æ�*��1Ba p���x3U��!� t�)IS�>#Ly�W�5׿.��m��D��N�8�h�=�[�S��A�#y-�B��p�j�+�����Zl�����Oµ)Z%j�����Q�k�YۓѲFo�+������40�1&[�J��5Dr�L�,;��Y.0�?B-d�]����������w��~̿���o�����[��:ʎQ�lܱ"���o^S��\�.Ї���G�����������v������M?� r�����Z	��H�C%�$���߬��j_rLyF�h[T"���8�����ȹ�ɋ=I)"ɣ��JM`+�v��#h�D��!b*���2t6o�'jQ�����0���U۬K�
r^H�2EB�,3�9OT5��	������j��ݴ�١z�!y"9��@J�_,�x��������d�q��!�=��mZ'��;�K%���*�U��#;�W�:ہ	�L �+��z��w � ,I���+j�1@UC@�@>����闷$�����h�mɕ���+�3������a���~�7t�p����vMl���i�"u2�1]v:��&��咽b�qXMF�e4@�(�N�%	8�;�bg;`�����������1=��G��z������;~���p~ZjD�2Gk���+
ZW˅^W�Ap���r���x�f��1=�K��I�7;0S��-yѯ��-��p#u��$X���������ufl^ބ�(�g�O�*N��s��5��Swx�b	Z��!ոҹu�T���fѾ�rO+��~%�����޿�-+�i1ǽ_:K/�N�5""y-2$�H!P5�/�)Ws	�Ag�<;�ڜ1�pu78�X,�3�x�ہ�7t�?6*�(j��.��a������Mh]�~�v�.�NFxs�j��]�vfS1�M�:�S����0M�	v`B��ӧDZ5�eகx>�4�(�/b�ұV��t���bʣ�8cO+�#�x��Jy����v��H��u�*=�WLk�D_y��r?Ւ�%sS�+q�j}W�qM��j�5dX���*�pNJ#];��@*�?Wׂ��9���$����ͣ��+O~e?�:+�u
������'%�!Kq�_C�Ք�&M�j��Y�o��MZԘriyﱞ����0X��)���@jF ׅ��R��\%�R�ow�PE���Rd�����K�Ǳ�:�6�
�䈴�)'뜗6
��Aj0xvQ����CZ�"f�,���Y��7��S-�y��ҙ�Mi�b�铊�yBVf�+����#�8`Y�ZR��h)�~�Ǣ���g~O����%r�>$�t��};e��q,r�,�MIV�nlx�-�4����R�3�,Q��>b[9�S��a��.��(�9�ۿ��/���qi�)�Hn�lz��+v��M
��e��ߋ� �5l���[k��:����o<:	$�C�����RL���:�"���G]|bƬ�V'�X4�ʎi""Y�B�՝Ƽ�h8�J�k_�)�w1�y�㠃��n�!2�"(E���@�U�B�8��k�4�!A¦+,1[~�>���#uX.IVv�±��i<*=A��}!Ca�@fJ�a^�,>��d*m+� �G�L"�0�}(�=J�j�>cP~Z7�U?�gn���ƴ�;m�pכ@K^�@��YԸ`��r�K���j\X��s�eB�瑰�����J�B�w~�[*���G�_RbK��͡n�%"� ��Y�k���ȞP*+4���P�3���u�7*ī���wF�?8�dy<gPcJ䉢���fط�uL�5:�o���~�.�.���&�II�';�2r)^���T)Ҥ~�b+����Oic��ѓK����ʦ{~���=���H/��Pňeh�>
%��H�)I9a4ޖp� <�b&/ ����'�=&l;���\���lTv�v�C�V�J/eu�ٚE���^O�iD3��!�Z�+-g���:U��_�u��k{3/�\�O��l|���m�	�i���4	���;4c�0%���sa��3���3 �ѕ�/kr{r��>�s>�V���7QsK]��3���W��2[{}vFGD���:g�?���p�֛�T���&V�H��.� 7z���w��5����^�9?�7�cJ+2S�h��?������t{��C��Ã����L�I[q	�-��N�TZ�����F� �?ٝ0��٪hףW����� �2`�9zMVX~�h �d��R�mP
y�lr�.�eܩ�II R��f�x�� {�T�T�Y\G8@XJ9@�v��^�Xէp���SVH�?�^Ί��zg��
`j!�}e��ř���\'Φ��Bs�SLٷ�����{W�����h:�vH.+o�NGei���ZK&�VBZ���0U:.��5��:x �i��w]�����>ࢦ��寲B#�|R�8P؋��]��z����Q��k򾒗�;��jcܬ��,��{b|��gDf��)��0;�g+Z����<�q�2{5��~lS8�,/Gr�a������a�äY��Ζ�jW���n�����_�i�Y�+z��m�[k�5���������]�R�,�^@;���0w�C���ֱ���SA(n�޷�� }��D52A6(z�y�3���mrT��U�S�e�3h�K������e$��X��j�(�sSѶc{̒A�vbx���\����5%LW�����C�cp�u%巀�}E�u��;�_v��`�&m�V�au#ԲH
�:_��!>�٥�❬c�X�I7u�X� c�tJ��
4V\'��L���b�j(�H0��AZ�o�8�	��]_r�!C*U�N5�K��������*��̼s~%~���	���n�'�25u>�j��$��a(�K����,3;�����w���d@�\o,Me⡔?��nϩ��U\����{���=�a���f�g�;'��mQ��9#���=J�94�y=QxQ�Q�ZS�<�Ծ^�Q�ɱ�ڬ=�u���FI�廳����Pjh�l���_D���m�	�?�B�~+�[X
za2?��2)��@5]z�� �^��Glai:��v��t'|����W%p\Z�:)�4-��+� �#��O���l�o��ښ���uU�U)�mA��i���Ƥ~�	��X���/]��dم-
�J1�,;�;��?!�t�|2<���=�y�ti-��V)����P�EX�i~��#k؃v���?Fv({��*<�z��%k2@���I��x��6�
L�R�/�:�-��A�D��)Ws�K� ���}��еWŪ�#����ơ���#b��j���v�V�8�o�B���9Z��:N�?��i=8tt��@�UP.���&&�(�0��a�u�î�v�$CzY��U�!#��xB��;Nk�')���@����ʉ�n��(U�(S ��<"��yq��m�KWC�Ƹ�[�C��b��!�4�����J)�1i���P?KXv�����b����h���G:@Q�%�}�:०�!�N ˣF<=fF!���;��$��`a�^4����>v�C_�?d�sTJ��:������%h��ԃ�o�#<
�����A�C3<�E؝�i��Y��ET��^|��������	��Y�A�aw���~�{��D����H?|L��%�kS�����.�O�V��ޭ q�=�S^"�<��ϷWT��3�/~c�H�k�|��C���ϋ��=5�MK��{i����j~�B����ѷ� m䙔��H��@�b���i��&����#.�e�]w{�p�5�&�s�%iP�GGt\;�QQ�j�
�L��<����+U����l�E�1���:����T�F8�a�&&*r�<�@���c�b�O/d�\�z��+���Lm���@3`��~^�[y�i���>�ff�K�ȨP���[��&_��]�:h�&�aЕ��f�Dj�P2ޟ��W�K�f�.�m1"�D?Kt��{+��	�������ZWӺ:@��θ��&~��cH[U�����k4rP�"�3Q���R�����k�'=���J�˥wWD�U>&+�LlL�+�.������/L����ɘ�Ğ(0���Gv���ݐ����r�bw��Ϯ�v+z5h<1�`�s�C�<W�"��yg]&� 6]�; |h~� m7�=F�����N|����hԗƘ��u��#� �*`�׽�o���~U�&E� J��t �V>;�|�(t���֢(#E�����0aME P�)�yZ��6.s���"����]iz�fў8�t<�-p׵�h%W�k�ń�������)^�B�y"�;�L�ģQ�)6�/ݓ��m�.�45�-cX�fQ6�mY��+�k�GG���,I�G�rI�FR4�_��k@��q��:7p�)o Z�*���ЇI����=yA��E�A�׾����ӚF�v������������F�/%�KY47�n{�s	�o�
 x`d�~ ��^��|�Mh��t�5 �Aߐ��[La�l���kV^k^MҊ��T�R\��_�������f��}H��Qt�ܴ9I3�=)k��<c2�=o��袵c��c���De,���;t�� 2�t�%Z�C��&��r5Yd(�	7� aX1>�n��%<?f6�3����=P翂'T3~ �}"q�1"�Km��21����l�ܑ?�s��������RT�l>IE�gk���ve��׌EH����-��2���YSws>H�:QM�m�*s�%�� ��LW$�>�&��;��;�Z��d2��AW�����l��A�i��\ii��}�d�6m�&��5[V�g�#Z�P(WH�rc�����Ը���a/��9�9��A���mo�UC���_b���R�s/�_�
}S��JS�	� �dK����_C����ZN�Ǽ��h��R:�`�z)=����#P��,ٲ�h�(�@�.i�y��>��;�oKB���W�;Z�,Fީ��{�m��� L�#GAe�m�PVS����$7Oǂ�AЧ���$��:̂h�<�[gU�/�H�#�[��!��k����O�N�H�;��Z>?ܾ����[~Ѷ0�{(�7^_��=���#�WdI���$��=���5r~
�N_~.$�0�B�V�1塘jÙ���I����B֒�N��L^"F�k�ac����*���@x��l^��d�C������6&�����֡��Q���ي��~��vC�;)��f<v�����|]� h5W�;�i�`��9@䭯�!2Db�o�C7g8� )H����ˈ�lp�!�f>>�i��zD}��$���@��,C��r�}�@���۝�����!p{e�Rae<��iTO���B!&�Vf�u�wl�I��,%����=�8蠗/:��]s�^�^xJ�X�)s]0��}6d2���]Тn޴�Cz:>���o ���h�k+���ݰ벆;&���~УLn����9PEf&�ܹI�m���!ܐ���J����.;����ɪ�@ޝ'�A{��v�E�ݴz�s�M�$Ge�װ����hJ-(+f	O��������5n.�`��F�E�T�j#�"�]_E�&��������C2��^V�3����<�B�M�fy�� �I��R����7�`\���*s0!,(uj
U��/-z\���I=GNh*m��i:���Π�x�Ǉ�9$<SI%i��>@�H�v�j���5��N��n����N�X����^����֒H����3�q�Y����_u�&~Jk�˷���dr��+/4��T/L�<_��ż���!�J����54�z�u�Ŏ�R���ڹ��ܘ]�tQ�٭��G5չN8Uw�Ĭ'���ٷ�=�����[HN�~��5s��[l:�m�Ex���ߧH�!In�j��I���j���o�XlxVHYEB    674c     5c0z��}�d0D�+`D��P9t�/�h��R�t�:�w�G �f�,��i�������(vGWDW��q��V�/(���a����V������s�X�Uz�ؐ�K���|z	�G�gw�(�I���$_�׀�z���˨8gx��9�)��7����aH|�`uQ�#-���4&�bpk|����4Ԑ
��|*6'��52q����ʽm��n����~˚=
�_��	�T�����sS���ۨP�a��[-�D�G�Ok���8~��41�xh��z��RM}�L��\�C���� ��p��o����Kk2����Ɉ��������* �jա�x����!��zL���C��Ī��1�s&�*� ѵ�w{��c܌p*%bG� rBW}Z\D�;�6v���'�>�D�gx.q�%�_E��=ZR��T��<%X-⑥I���~4)��_�gR޳z��� W��):1\�l�v�?!n��Yc�/7f#�KS��2z�9Xo�4Q�X�¹�:���� 7\�G�V4ݯЙ���I����,���Z�_���٣M�}U�;@��0�B=�&O_�8񌲉���:A>�״��E�P.f�^(mV�3$�r0�~��O��{��[MVF���=�U(�I��@w���h�&�IJ�X��uS�~}�+��w�mgY���Y�s��ځ�l� �,"s����Ls��%.����_�N��ߪ�;K�ͺ\p�Q�jڃ[*�w�Q����:�������)v��cz���t���>Ŋ��l$�^Bۚ�S8��� �@E��Hq�Zi9y� ���9����"k��xU<�/�Q��p�	��A7����W��u��%����2d������n�3Li�C��7���ƺ��O�M���3�Μ�Yq��V��p�c���-b���1�>>��<�N�
��Θ"�X�C�O�ֲU6`R��;Y�h-���z疘C8µ�ԏx�M�(
�ݩΫ���0/:G#�R�B�J<-o��1�y5�����7vx�WҦu�b�v��7.�@o[�\��.u�^�v�,c�d8=|o�l��	�Ie�V?+}JRY�7)�R=Y�[;�m_p"PED:<�z���nu !����f��d��N347���;�iS�ɮ���_�"ϲA�u�tGP9��I�)b+����G��mK����S {L%ăB,�8%���t�W��D ������ް�:B�4��7\���/Y��@��[��O���]�ȉY��:��|	�������ܑ�G�b�}C�obbh+���֗v�;���B-��~�*>�����Z�C�񄗼�vb��V�����38�u�"R��]�*`
���e��E��|K:~qiɈ�{���n\Q���̇�$I�%`�O5'����olO�M��z3
��$̂d B:48��R���ql*<�a�#�T�w'���V����$�