XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S�n��(�]�����`�aa̦�3����)��#=�а.����#�>�3�M�A�]��ʖ&�|@��_^�|R����9^��ky��|�eӱe���BBP�XZ�"���"��%�=EG��w��Ӈ�e�%�%2+#����ֽ�ރ�\2�?��|H?��-C]d��H��U'd��,+)�{X��4��l�S���Dfi���G������=�e���>c�!j����Ҕ���i��X��o����1V��2�G{��f����=��v[u����y�/���p�$���5���^��u���w"P�tPƀ3��,���(q�����P]Ґ{ o8������'�uC��YU�* ̃��AP���G]�A����i!�&�fL�A��\��
�l'9[�n6�w��J�J�J?݅��:��y�����j��Q2�9�W���w�B_"~��ڔ����$�����{f�`�?�
�X��vT�C�<q�;c�À1&8ߋ��`�a{I�v�T,���������%d񛌦�t���[7�N�6����|���W.�Ue��e=�$�k=�[�0�7���B��mޠ�V��8h?�nO9a����ZO���ל�mӪ>�0�Td�8<��1,dXZ���R0:R�z�RkKi��'_:*������t!���kj�s�D�`̛��n�,�G˄y��bj��6��K"��yhB�8�eT�s�%�������D���'��i��&��+�<��7+�D���M�&C�XlxVHYEB    29da     af0���p�z�6��fc�kN/���ҽ�6���W��~�jO��:�*T��jbؒ����Єښ>w]x���>}�P��v���Ra�g=���H��)�[X��L��ܡG�?�+rZ��Rtzv�r�Nִ�%��c�wt��2K,	Bq� �+�g:���W�E�)خlMr:�Y#�=�}$��2[Ժ��̬����8�?���`�#���Z�Nٓ�y$��P��7y����B_.l>�����C����|%�fQ?��ޞu�~�X���'�tR=�ٕ�ń�n*$�m]2�����S��%>[3�9�,�}��i\Cѹ3cI�i�er;�jzA�ɦl33�س�Ω}5��e&�j�-n��@���R����Ϟ��t�c'��g�_n���.����sI�s�}l���(��!̽�\� 6��6������A��Ȓ�w�I��z�q ���F��|���6�C�f����4��8ZoD���{{����D�����A��A�^_��f�0���Qg�q,�Fn�vq�GT�0N��� �;s���5m7��`��<W�8�m���AV#�}������Wd���T����g�Z1ej
%����Y4���p[	,Q��G�������D�ظ�	��ա֦Ҡ�wB�q|�[��|��cا���-�Uiͺ���ϗ��w�e���doP���_0��^�
�|���~&��~ץ�z�>g��!��IR"�)T��Z�Kap^�ڣY���p8@Ιhv����JkZ������?�i󚑚�ƻ��Рٽyn{�2[��ێ��Bz-5�=�5-�E	h>��2��~L��Y`� W��e�U]?̙b����;�ԥ�0� ���Ȼ�uQ���m�O�::���˹�\��~�mݛh(��hf@��e頝i���<@�5,���B�m���vg��A���5�k��S�1�;«��4��1g׌+�W!��FoW���O�(�xE2b��O��ue�����J�{*me�)M0�+{I�o����+`ur$CYI���850��.[�O�,�x�|�k�e��\܊�de����2N t|����Z�Ĝ(�Ķj�w�1��)�(��˘�^a0��v��=�2=�g_}�F�{�&��0�n��}���=0I�a�X�^�+V�럼ϱ��X@��j,�&�h���}�o�SWNA�Q���?Ω�d��a�'�1(�%��|E��֙��n��sL�?�+V�x�wϨ|���B�&�[�
�� ��,(���MV����H�	i��̅��!Umҏ�����)I9*�R� ��;�ؕgC�I�B��. sq���6���p����X�^1s�'9�,��0bǤ�`��vhϸ"Z;aL����l��҂JU>�Z^�Ov��[��v�cJ���/��ι�y�t�S�Pn.��U�ph�������C�%��r��%�&PY���<#�_��5�je~�,�=<�i��%Q�Թ�Q�
SL�s�.f�
t�^JeF�O�m�b+gv߄�3U	�H��/��_�Yĭ�ϟ�"-jR����'��6O���W��+<`Z�]�4�#�����~(N�~ʐ1f7��!@�A�t�w
��7N���Z5�0�K��]u9��
L�z�ր�Y �m
��������(�y����ܞ������ڞX�%`s�M�BC4��r�ie��*8�{��K���,A9���_+�3��ժ�7z�w�E-ṩP�'4��T��9�����ܳ7\Jc�N�0��)�B���x$g�`#�~�)ۼ���]�c���4ޝZи)P4Y���,�������FAP ��)����{~�Y�hu��;Hѻ��u'7r��[Bok>Y�8R��u&�i����R�i��-䫮�&����1U�wn��La0t���'Zz�O�&D��j���=LKy�D�	�x�wmA����Te��-Y��!��-t�x'}��ץ����6�����[��@�e�;����sz��oM���֢�\�8¿Hw���Y
Ţ[dF���8�#��
�;1��WC��}�^�r����m��K]˽4��0j1�w!�3�� ���V�\)aCr�����F���m�(���n��#�Ś6�ej`2q�mթ{���Z`�"�m|���$�u�>��qZ�ƛ��}'��\>��A��T2O7�u~*S��\i�/���$o���ͅL��ž.Ft���k������1 z�L�?��Q��I���~�ǔ�>w܃{d�t�������C�Y����\4�һy��a+�т���n��{ߧU9�3j8�B�֪�K����C�ݖ��(��p�.�w�7V4��UJM�x��!v��~21�g��CVB����y:��ɫ��Q�''����}>�/_~?y�d"~�~׶���z�D�g���������E�M�C�.��)����kӎ4�p[@j	��}=��j:P(��e�Ob5��6�P�R$8�]�t.R-�W�L���:�5O����jjϞ#Qg���$���^�V���f�'#�o{�C� bAC��Ћ�!�-?�Qa�O�>�YԮ�m�콊W|����iT�bX��Δ��t�m��� ��x��o&���� �����=�o���/�z�;.O��W��#2�%���6r��f.�U��1Jw����*�t�h��S
�r����?qi#a�G{�U�V�~D�ӵN9�j����F�;��Uo�pQ9���R�÷8��N�